��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�)	�ŀ)v�ޑ"^��F��L�> Ó�����M4G�h�.Yv~��f�+�E�9�?���;�Ω0�4��H�;uS%."q��Zd�/�]�+G|��Ԇբ�n�<!�?�a,��5_��=�n�����~t��^}��ٸ�/��eLУvi�i���m�ޮ%G����i�}	�71\&��cq����+�zE��<�`\�L^�e�|�ی�k��=OV�B�v�@�1�^'盾�R��9��'E�򛚤�p�E^΂�Ok��������aG|#�	[m���}�����R��=��ئ4�r-����[�}�x� �|�LW!�c\j��:���ȳ�oi����_v����jqQ�#�d^��Fџ��<0�
)ߪw�B��ֺo\�s)��M�[��	�h_*9o��E_���]��F~�#?ٌp�&�5d1�)G+��� �n���?z!H��x8��U2�#��#T�I�%j=�մ� �Q��9n��C�)��Y���h2�'����lw��9\7�� �9�`�ꌗe��c^E���2;�%�R��� �w�Pk����9���sr~P����u|&��S�-�}	%N��v��	T)%O̘z#i!_ ���*�w�3�Ļ4�L�~�Ǌ���R�o��%!��V��R�����	+ښu�u��a� b� �$ɓ���������G��*�N�
?A}��02��߫w�<s�O������!&v��šc�lA��&���h�"@$��H��r�l�f)��b8�ۘ7c ���|�(<�1��Yh������*�㋽.L��E0pa'E���d�0E�J���G�?�X��$�fxo�#5�P}����,����w��g�VN�V
�#HȎ��U���̏��;Y��c4�p�C��Y9�\v	�5�MX��Ǌ��%�1��9x��X���Zk���j2 �5)e�-oO�P�]�ѐ��n���F�T����
)�@�s��t�P�܆�,\F�Ehi1�������"W�_e�y�ͦ�>>~�/��};�Ӈ�1�GҢ�m�����
 \ n���&��z��e��� ԺU��欀�Iv�.��r�*����,̵4�E�,!>�J���p�֛K	����
X��^��/�YԻʏ���7%�e��)��o�nj����������w7��y��܄��D�s��ﹰ���n�L�T��۞�r�(�����$	
p�q� ��,��Lí�����U�4B9�9'n� 袾��R��ui�-kv*��%�=6þQO��6p�J�y���:>wꀰt�ߦPH�Z�f¢'��;?�ܒ�A&�ƚ�n����ʹ��4��.k���K��V2q�7��NU��"���j��o=C�����$H�Yr�G�)q�����x�1�*z�~(^L��#A��|/�N@�3ڀ|�d_or�vљh�b��|���D�����7:n>c�V��^��K��N��plx�J�اP�ek�[ ��)^���Q<D}��o�0`CI_�"c�����Omd�O�i8ɸN��c�fDA��i)�>c�/����|���w��4�}��8dx�$���j��h|�����#�����B��a��e������EZG3!·<����vf#.W�]��n?�P�ti}������]��~��e�A%8}`���.Y�V^�OF#��>3���&&��6���.WbКp��p�ڊ�0�FT�oE��=����8�Ng�uf�L�*e�����M���?�vЙ��E��Uˏ�X�.���a"�x,pE���Ak~	��������e����
$W;_�S���+dsy�%S����Jd�	[e�9����M�D;hD��n�����	�ճJ�r~M����~k�s� ���
��� �ӱ,u���l�|=F�$f��b�}����������2zU��2 
��]x�ޔPM�7��s�d�����nl� ��{��yBv��m���DD�Њ��?h��F�E�C���vRAH8�to��s\�s[���!�!�*4�u�k�dai�*�7��7�HgLȧ�4���B���Wɧ�s�0�T��gS8�綕0��U��:��[@���0TV��R��	���[���d��>W��v������h.-K�!i� DN��aZT��q4a%�5V�޽#B ^��QN�H�7�%�Dc���R?�)Q{2�!m�P��{�:p���xR���,����{ �s�u�a�_o��m�ssA�g�����-	�ҲB�qC��'N��2�6�[��9��Co5�r۵�ں�90��L�_�6)L�;jF5P�J�Ɔ��@��X ����`�Y��zt�<��tk�����2����nN+�M|Lm��
�	��)�0j�iXKd^��k�~�~=�	��;���(�H��)fL
�DCw��Q�
������4��-2��.,�`�O���������X���gK|p�SX��y5�)����G2�z�֩Q���s!�|.Y�P�:<��gȍ�}¯/��5k+W��&F�A]�F.�9 ��6�Z��&?"+����,#���uҊ����`���a&iUo}��:qV#jxQf+�ۖFwS��Zd=���rdy�h�J�:g^Μkbs�BK��/�,/	]��WE���&�{�b~��3T���e�R4W�hA�#�wН���ʸ�90V�M�K��E@l� E�KF��Q�c���l��j�1:�����D�Co��:����y�
&Pd�����D���AӼ��m9��Ja�q�+D�)ƺ��$Q�e-��v��
�L��M�f���J�.�B��O��*<�V/ �_5�ܭ��d�XH`���S�a����h;�j����K2������KkM۟m�'{w"��y�1�Wz��G���/���.s����lK?�������n��8���v�	��G��pva�uw����In���!�Q�9��J��l���o��(�}°��K,��q�L�lE�b��֢Fm�r�v�t����x�zG���buC�T�Ί��n��4-�������[#�H��fcS%�\&x�c8)o�m������d �q�4���F�7󂩡p�u�'��l��ca=�Ip�v�4��׆�����&��fW��EG��_�3����m�5�Ⱥ���d�J*�'U�� ���ƛ�Ʒ=�w���.>�������xI�4���	[w�0����l����
@�d��H9 ��C�vC��X���RS����k��:4Vx���,�d%N�|p�.���7�J��o}�8+ϱ%�P\u`���zU��(7�$�m�&���3�e��O�����u�6�0��{�O���MR6z�?5S	x���W=�n�_Fqp��@���8�V㓴zi$>C�>��J�v��β,��vZ�=��1,������
�Lk#6�\o�DS<�(��U�GQ
�u7p���D�<�)�Nh�W�I�a�W��/3P��[d^�	%SJrQw�\i��Χ���
�����ww���+3�� O��78��6��3���]R���{�PmyW�3�m���)����'�Bp�J�Z�3�W��A<���HAAT�{�)�^j�r�o�o;�p���D�z���
ƌOq���H���0:)��+M�G���uz�hg�P�ZN��\��������7Y�.p\v!~ݔ��b���$�b+أ)gd�2~d����4���RVH+�vD������Z7�w���ekr16��ɻ��6Z�0��� 7��d�:߻F��l<P�%_ �C)�9���߲�ʅ}����}��v�6��%|C;<P��K���Q[C��mҤgb������Y;�N�/��
�5kfDhHL�1ͥ=�<$4b��+<��I?�D���-���y��rO@x��y��䩩�{V�;��S�/Op���9��ϡGY���я�����2-�X�%�uEq1RC%0�/��5�%h��R��Us�l,��V3��ʖV�#�k����U��ܼ���
=�U��>������^��NM3�O���ɶ���B�v>@SN���Ht���k���Sq�If��v��"%�Gꡅf2�)�:��k}��v^|4�`[w|LnB����'��-K0��������$��J�����Hj�lpfG*�5m T9GP�ln���Kޮ�^�I�d�J*�ڲ B�I���&���K�	:s�����sj�^�S/�(P>�),.?QA�sNo��.cz�����3��az::C�}�|����O�?'�Vw6{2�[��b�����F�4ߤ��b���0ƪ~VH؄J�ʖHm��S,u�I���ԍ�i�asq U� 	�����T��Y�5w��l��dl�1�-j�qw7b[9Iw��Jz���Ag��؁�$)EX���� q��ؽ	�����N�/��-;��~�:���ڸ;�w&7j6�߅��3'
���TB�?4�j�UjM8��Q��o�^���(���0�J'Q!�}:�X�6�����56-5-���^���d��>@��%.�<�\H��nZVFx��/N�BN�~c���?Ak1�Q�豩>��ţ����33B��Y�m�f��b�W�6�Z�Hv�:���ȉ�1C{�-�BEw���I���:Ĳx��*�<]�ݱy��s�Q�7C4u����$nȞ�".�1}EYA�I^�ȵ�vՎ�Y��
x(>e�\�H�����3P���p�wCX�J����� �]�����4��E��t	kx���� ��!��9��`V�)9�[�q�6A�����^�@����d�����U�#�i�W�*'[�կ�-��㲀�.3���ԯ�5�%������KI?��N믮2���T~�t�� 9�j�n\����%��`����SA�:V�1I�1�����!!��m�oБ� $��[B����F�r$jf�K�(���s����Xs��[s��A��	Z�*�8�~��ހf��R�*��G���n�H�y�*��O���93u��TuI�~��&�q��lȄ��4eG-��kʰ;���N.�Y2�묰N/#�+6r��IY��p/���3�}��B�
�cl�;�8��v��i@9uR̃/i���*R�]&h�YY<�zo/��֫X#�Vس:���N���8l��e�ۤ�:"牎ԲpI9�AY��u6�X]�%<C*�+����RN�Z�#w���)k�T�L��'�0���)��;�2���l�4SL���
H�ӂ��BZ����]^YI���L}����4f���s��|jH�gP-T�	ݓ��^\��o��G:�<հ�X��T���'7�"Q5d�ӊ�]IBĵ	!����vy��_�wg�F�e4[�c+�"rrCV�0������Q�Jh!��}߄�_���WP,�U�CQ�LY6��n?�%��9~��F�SG�>����?�ʰ�a�:ʠ�º.����i��$�u��a[���r�8g�ܳ|{뢸5_��_��Jjbʣg9Q݌d=��1�˕�5f.��S*�������:(QՑ1K�(k��dxeT�s��v鲔O����vQju��!;���R�Ő&��Yz���"�8�A:��������������_Y@*L[ T
�Ru�<Q���j3���7p�ݟ߳���o�p�`zIu}��.�3m�� ��|��+�B�u�����&p�d͐�!^����T �GS=�u�j�B��Y�*7���}��T���k��ZtpO�3���Tl�p���b�^nwȪW�Y�`�U���V
s9c ���'Li�S��������KvlK��;+ ��n1U����`T��T߽�tw�sKl-���J��������ҡ�6�G '+���">i�䵠��YS[�fmo�#��4��K%��.��ײN��j�)��M--��)4��!Pс�tc�iv�t�������1��k��H��{�N�J�S���h悃��F̌J�:e]k��b2�֜�_r����V2����o̼�EBOr�*Zcރk�>���'�=�l����@3��{���>C��vwn>���X���X�D#�o��Yi�<��ҥ��5�X��&c[�fR��A2ԃ�N©��4yO�Y�{���Ǩ�P`t��pz�n6���� �>�fl�#�k�Ko����U\9�N�#G���hu'L�X�r�[j�QM?��s�L���u�OrE:��sO�#�4�Q����� �ڵ[b���Y����^�L��b�t;�!_Y��I���$���	?�0�QF�&J�Bc��K�,�4y2��F")'�ɢqD�D�5�\���V����Ьb��/�%��,xpŢz9��9#b*����D�����9E7������W���Ó����78b�߿�s��x���2��7\q��9���5�h�*.{��5u���ڹ�n�r�k�A�\[��c� ��M���>Ӏ��F�&�G�;�{T�����}�2�{-3l<�<sx$~ǩr]l��]t�V� 6��=r	(�n�P�2��}o��>��L3��I��?��o	�w���K���`����3���JU������A�49��ں;��g�Wf<�i��ޑ��@�D�-�iJa�J�<b�@(Cd�?�C�U�����2�c��C���@)��L�Q�yb�I��@�Ċ�8���}$ӉI�=T_�����ۭ$���K��#KD^��5�j�hfTW�=3)+��iA:��:5�����ʁ��Gq:ʑ���(������+,p#��Em���^ؤ���3Ig5�Yr��dU�����^vA�ٙ��cs$ى��幫#�WgԎ�	���F�[֣���U�ul|P����xU�~R$���:́��Ƥ'Mmw��=�if��-U�A)�Q�h�pz'���hEȭ0�в�`eGE=�5��!�ux-<C�r����PJ�{i��n
����*c龼x
�]����R�d�@"&1�5��ګ&&q�\[0�O,h<�,Y�dA��m���04)��՞�/�m4�'��j��sE�V`.����:�Y��\` _���$C�j�۩,Ef��1�=�����#�	!X���-4���˶B-�>X/�L�`�fc�vvv<��Q �~ý��ϐ��vU�A�OA�m��� �;+�(7zx|YK�xT[� 4�xY]�<�)���KJp-���o�.�i���?��`�T]�4D�rjl#u�Py���:���`,�'hR7��̸2��K�	��@�fED|���1�8aQ-&�{�#�6m�H�v��L`B�֠ݚ��߷ò'��W[�
7
�}�ee�t�H3�c��qgBi��丗����tV~0���[�������m�J3x���z�H_�d���%�<�.����������F/� �u�.�z��9�NC���)�[��3_Ez?=�����I7��66}��κ-9A{���E����r�풗�\P�\���4��U��.Id����s�Bf0b��|�NC���`������;��ah��Mvw��~���p�2���y_z(��(�e^3ޱ��^dZP�7���C�,���x��� ����Lu���,�gb<퐔ϯ��jVj1����U��ÍhÎ�L�w�8�*mt�V�@[��(����/�'܀���.�!L5�8����'08�X��.�h
��V�8gG���:,���7� ��/5�Ǿ-6.qZ2�`�M <������O?_`��XND��|��n�+��
��IF��f%GF��jgV�k�����W�9n}�_�Ѫ��604���qh� ��8ŜeA�'�~1Ol�+z��jЁ=Pn5$�6Fk��ixO v��wo\�Ή[E�t����Z�˻\�3��Ov�����|��>�28�	�gP�ֻs@P��u9p�vk���Y��1j�ѓ#R	v7ګc�ӻG�[;QW_���1MHC����Y�n���n��3�������L�X燤&y��)�&��^�=����*�с5���/�[%(/-3���89��D��(J�{��5�l��w��ɤ�����$�j��:��L3��9ȈCα{��7�0�B���KDR��L,��_�˰߼M���69�y��Rb�T���m8�eť���E�c�Јk���_���R��dG�}����*N��Z�KA��O8Z���%�����i��r�w��/�U+�2�^?��c̹N?�Ҵ>�)~�1<9}zH����S>�s�'Z�8�X`�6 ���+Ϋ�8x�EzL>MO6�=�t�f�}�����87x��۠�ρ(�Y;M�k�Yj�����xB9��Y�����4�K~��PY'���P���S�p� ��8��]���[�$J@����0R$|� �YN��"]ݾ1��19ئQ��#b3j��+L�.6ǹc�&I�"k~|@�-ʚw��e�j#�����Q�4<����k(n� �.C�6�>�f�H�����_[��.c�e���������aH��g�S�W���r.�0gɂ ��8�gi��V�������޵�?�L�,�3f�Q��(����tP�hpp�p��) ��_c�ȱ�9ʵ �ʄb��d��1Hͪ�hG2�3Rr.E/OT�w7Gz�6�������$�eZ=\jޞ�٣ �Y[�0	#x�K:����m[v�3��N0�D�؜c
��G���?� m���CJv��a(���3-nĜ��L�׀Žю�G���i���o0$y�FP��:d$� U�y�}�l��2:Ս���7��a�ޖ��#,���o�I!{	mƄL��C,j��0���5/:n"6�:������l�Wn.ݫ�:��I��&*�?jz�\M��A锷�J�|���&I�D'AKa.�&{�&�0R��>u�?&����W��z+6��$̮��[دa Ɔ+U�A�z�`�?�Xm�ȫa6ؑ3����"�WT���~b2M��A0d#�0���O�!v\x��VK� �N�se�3�6Z���2Ӥ��$���)F�e"�҂�6B��$ھ���/�
��=2�HW���D@D�K���W��fq=�d�M����&�I8�u��Ԙﾫ�����N�*Q ���W��4�테67�{�x70p��I�dIȼZ�n��蔚T��R��I�c� ��L�/Z'��YF�gM<(t3��	 ���1]�P�����]��ߤ��V��5�nz����f���r�2�����tx��3>�u/.�7�tT<��\��A67�;�u�o�ZhS�%DRg/{oy�#�[�eh�jBI��^�5���7�$	'�DJ�x6´�G5H���h���+�!J�Q�a�W5�(�&��#��	ȍ��C��q�� *O���%�ؾ�b-�?�L�{k���ę$i��3�-6J�S,�֌���?��DJ���4=�Q.��;�[�NpW��� �yՇt��-x<_���x��{"d�a"���	�a��=��0!�G[��qO��-��`��Ҭw�8��X"���2Ƚ��%�v��0��{�!"���埑hQ��X�~'�(1h#k�Y��7�b�
�u�+��H��]�R-%�aE{�ii�,j�ʏ�2���|#v������TG�))
�y�m�p���9���,��i#yN���a��1�� ������*�f�iR��g��F�w$�/D焝�Bt|���K�e�ز��jE���DɈ}T�#Ԏ(��E��lud��%���2o:���*��D� �E���l�X��o�u�榷㦶�yy��!��������F5������_�o�tJ0�wǄ��x���y��4� 4�=O4�VR}�t�g񚩔[ؘ�.��H+�kw\}�H��{�P�$��I�1w��x�@�K��I��'�N��l�JD��J��$��.Ԟ�r��}_����׭R��@�9|�zJ`!>����*[Tb�[�7����|���/?�$�k�^��9���n�Jl*}9���'�`ݸS8�T�"�V��i��9��2JOx*����{��T�E�v�4�R4�bX�!�	��O�	�CO,/oe>��Jb��d�$Mf��e�;諈څ����(7u��uUvhq�������G������ ��
ٍ�:�Lyȶg��?�-�W/d@vuq�đ����V�3�Y_�d�5�QR��/�'���}D����$���E�,2k�g-���D��2�N��~�����E^�hK;~G�����!r��V�E��C�_>�����{���y�<l���6
&>��sM��=H�[� pM��$�F�(]����U��x�ĪE��
2��S�""d.q5��$�،���B �h�BL�Ʋ�D�v�$J�5\�b����6#J�e��U��{x�S�A{l�\�>[�K��g�Z���_���h��	֟�er�!����ۻ8hSh�0���5� �2��$%��5r#�2��{�B#�ĳ�	 ��5D�
ބ��&�P�l��qT��KI�,%��=5��&fI�w��I���B����P��:�">x.N�?�>�G�UE�:�=ϷM.�F�OM^/���J;��q�ٛ4g�
�T���8��l�>�J*�����]�`-���8k���/�w#rV;�+ѷk�J��s���%Z���W�=�)�C�D��TGE�#W��lHN�G��:��ڷ��P>������mQ�������/������A��6�{��|�J�ŀ��q�a�qH�����
�5�\��dc`�r��u0�*(�'�U�΋�9V������Ċ���Z��",�u��0���nx�h��E� ��uf,:1��x1򮏅8B�l��#�~}

�o�)��큰/���#�&-v�*��Xaz z����x�r�J�4Q$��U_��*v�O��.�g��X_/9�Y@C�z7Q�0��� �HV�C��KME��+�O�n �t�K���j䩫����xUⓦ�����p��s�R��d��9��v�&sew!����j����K8u�0�:o�����ǡi�u끥�~���[�9��mS�˵�����`���Қ�_��~��.u~�G�WK��1⽞��_�9�V�8Xt=r�0�n�� >?��H�ۤ��u�_�̰��q�q�����)Q2�^L�_�-n��_W��	��Q�?�)Ya�[��/�g�}�48TmĴ�m�j#�hF���/���QX�p_RQ�=_&�V�Pg�R�5߆U?�k�@�T'�b��#�pB�UN<^����Ɣ[z<��n��3�l�z)����M&���9�Q]�w�;�(�I�?�G+�6�+Ա%-D�����q������M0	���!(���b[}�AX�ݔz��CG\���0ef� �o���3AY;�O������9cV �0Ghs���3:��F)���	'K@�-BC�լ�yS�������F����x�Z����&T߆_�$?]�xawŤB����ue��fX��� �S��u:�)�jr�Թ��w��Jd!�ػ��}Dx0���_�~�"t(F�"����.�w�DB��Qp\���&���ۜlbL��I��$�E��������������_�n@����n����p��C���:��O�ֽ_��c�aNS�Lz���!HVa�i��v���5����C�NK�Բ��N%%Qİ���2��/��6�M��H�9o�w��o�3�g�SE��T[�P�#����Kɪ��n&��<e��Q
X�<����̏h���A�h�WnV�V�Y��T�݋5:UG�X�!?�.�����5���xUŶ>��@8���j �j��zc����k���I�&��?w�2���
4!T�v �ep���l�h��ҀՔgf��ڪ���[��{H��g�Y�t2(Վ`qU�`�|�I����Wح	�v�*<��	�B-�d���׵��M�k���k�,5'*Y9֓�Uj�K7����z�����p�U�sZBq4!C8�R�ۃe�\��c�P��v6I�q�)���P�w��(�F�OT� &f���*�����.����tc�BQG���ڴ#E7��q�;ǋ?�+i*z��V�6ϱtx�3������v����&��'W�B�`��uW��	�E.�!*5[X�(�����/�>Q���ɴ�7bl��q��C��i=4�7�MKމ�������0F�h�nֆ���bv&�/V��Z�]"���~U�6 l{��G��pF��FE��{����p��.��r0\�
���S�����ݠb�wF�����3n�5Ԉ1y��]����ϑ!>���)O*]J]�H �C��f���Y�M�瑯S���6���&�)	�U�p,�zj=�ړZé
��q������ġ�|}H��E�Gd���&ݔ�xֳ�ų��	�o�h5����h`3;vCӗ�h���mG�}��"3i��n���Ax�`A��bt	H"	z�>��,J1�!2v�nI�P��D(�n>ؽ��F#>nZH��_�)�]ӑ��,\�͹LY�(�Z�I����^T#��Z�;Q���@�0IU�i����b
��0��p�˫~�������5����r�����K�Vj��`1D'KU	�����Ȃ��PqG�α�������ш��x����M�2B����{�Z ķ4�5�4�j� \˟�9�C���]�|¦��'��:��
��[����X��V=����4ufhN�&"�J�I#?T5����J:Qu��֘9p����<>,Z��v!�	"Ũ��W���Y%���!�����1;.��־O��Qb�cw^���Ec���G�{��\i`�Kk����o���yN���?���d�8�"� �f���j�vrq�v0�p]��˻;���Y��u�S�������	+Z�Χ�.ƽ��u<����A�j�~���}RQV����-��f���~;�>f8v��!j��+ܘ��W2�C0)����6��C
�4r�k��Ye$'��,T�Y��e�Ps�N�˪?!D������p���1�9�o��&%0`�}kW�{U��a�~#X"u$tF�7���+��Sl��y/�\��d���Oϋ�Y�S��_ZZ��;�g)���c3�:."[�d�Z�D��HT[>�bq��?��d���/��4�:�EڕL��VT�*�^�B��-��a�z
> �)�~�UXa�%?VZJ��������l<�R������}��6>�-�rr���(y|�P�s'��룴�W"�v�2��FM�:	�G>p�)�Ѓ��JJ�Ha�A�tI��є�g���i	��G��&���p�V!����h�Y �F�G��Niw�~H�3(dۚs</���s��NT��<���!9K:�_ă2O&�VĴ�ƟIg�W���2���9�Z��	J�����q�-��h'��Q��\�0	�+�y�L����zY:�@۔�S���� ��$aUt"�(N
��v�ݡ�KOwq�TG�l���O��"��|��=��Ƌ�~��<=
f�U2)�kc	�eJ3� ��:�C�7m")��]�r;'��$X�,�����Z��üD������(}��b�e�⁐A�.wȡd�Ƴx�
6C�RU�rU�(Z�Sx�X���&���<����ټ�A�.H��O�2a� =�/W���BA̚ڏ�vc��U�ì|�h��vN��y�+kv������.[�`�e�:. $��O�V����.�cQ A���y����H#�����u��MU��gȲ�d���(�W�<�W�g�/:M��	/��ҍ_������,�{~�_;-��+:U)S�wg�`B�ȑS�2��k������9���fU
�Є?/�3���p���{~�R����=?�@��W���c�k1�VBZ������6���6=�Tk��Q�;�|�͟��{*�#�A)��/��+�!�#��|k������[�XM%t�a��9�����N~�>���y�F��E$�����7M5�tŁ�����l�9�Y �6�T���)V�R>u���A���%cS���gݯP�R��Z��L&(��02c;5T�;A�-
2�h'�:��BGBY��l�|�(�k��˙��p}������Vz)t׬���2���}DZ�=�lm��G�8w�x1��=g�*�f����i��h��gcw��C'��~yS�����R�`&zD'[F��d�����U>�N���ʋ�� >�)�qa�-BR�<{�9x&��ܰe��(
 ]Z�9Qq˰� �ȃ�x6��v�w ������ �Si0���������'��F<��huh�s��o@Ћ�Ƨ.^h�>�+������o�'TWP��\�i0�1��������a�J,�A�0!�z�����az�[;D�^M�Ym�Q��p��z��!6�X��K�a)��� ��LU��ux�˙���>�B`l�|���:�*�����c	]z�B�eq�z^n�u5��R
y���'���'\2n��J(�U��Y��z{�M~	�����β
��3r02[�(1�۩Ĭ�.�X��t��Q���7���T)Է���S����Z��h��*�͌�]����Us�E�E��H�����MG�³���,F��V�D�p!�	�v��w<�e�IP����푋���3J�H�lA��S|~�6z�*�~�=��ǯ��>�X�	'�(��kbd���5����X��B[���p0����l��GQ��Xl���Kj۞��`�ڈ0�9͚��y�[���؍:knD���e� �>+��Z
T��{�����fa���U�\r����(iq��x���o��8p#���πT]��tQ˿4�b~�\��l�n`}xݵ�
�����d�崜�M%�t�S��n�&�@h������!�o�i�m�,���"N��EX��;�}���7[�
��D�;L6�4���P.�M�"��ov㰽94o6�2tn� o,sj>�F.z��s�����+`�HvȊ��-�H�7��髀@��W^j��\�@�.�qX��y�_�H�ygHZ�,P�t
R���ܯ���pb#ue����Ɏc�dء�]>"[�[0Ԫ�F9�`k9��+)x7�;������ E��R.Ӧ��jF��K��}^�%�i�X���w�p?�y���+<�g}�����I�z$�	V�I�Qo�$-U�>EOdԩ�"���;��ÿ4����A�\?ZxH\���u)�'���zٺ����
,�H.��օ-��/�A8:)�5������bW��?�Z�F�=���t����n��І�¤|.���\:Ծ�ƶc_��R`t^�f/L�����R���-N0�P͓�RV�Y�� `����?H5�5�-$c�v�"��k�c������X9�B>ݡ�|��
jQ2��d�M�iM���f� ���Jxw���09�`�s�� ���^	�08/a�HV�$1L�`~�9��FOSN�v>c�2X�;����\�(>1�%(%�,t�����A6����z�s+�_U+��Z�>�/@��H���:LNF[a�%w���#�ƃ\7�d`QvEpY~k+�ھuTwϗ� \L�� �������O�e�߱���=�6{H�=�8n�����~R�l�b��<�ᐊ�+��o���~i�q�&�"�΋��8k��J�0�p��rG�΂gS^V*���U��0��8@��hq�yi+��͸�n���F�+��4Cm�q`i�Ûɽ�ܥ?�r����y��%��ݚ�qk|kZ�Za]���;�o��>��ғ !�r�F��p
i=YOM7f���ؚ愾���N�a)����}�#�%f\�ˑ�� ��/A�be�t�9���N�s� �+��cm|�Q3Ř��jn��W�SF�1�T-Wexx�B4���?����r���_��W�����n��XT�2`�WgK��R}M1��5)���=PZc[(�q���ҏ��Ƈ���_,B22_y����
��e8j��R�	�k�q��\�8Xi@�vt�J� �0�D�yP���>���Q~���A�,:E۔S>:ȭ�>�@Ʈx�y4�¤r�N�5�
^��+@I 4��
Um �-7�nbx?ގ��X���C����d�ϪG�ܧ^��?� }SV�&�D{��/� s����q������_�l�t�&aO�$��� �r���$ӼC>�x쾐cM�p�>�{=�9m��:�]�rH���V�U��>a �2���&c	e�Ͽ!�.e,j�_���A)�SU�������X���Dm�O��BEx�ܡ�R��q�%h0U}E�^�ɱ��h�?�y�z���o[\���L�<����6����XC��gy�����CxW��Ja��E��ȉ����0���,w�ڍӐ�4�ZL�T�ڍ|h�׿����畘C�PE1YN�xh�:f^�C¦�.�0���t XW�"�;���������\,��G�^�ސ��^�˜4:��c�����rb	�`[z��#�u7e3�HMl�	$&N���w��JCT�y���N�J1�컬��c�ˣ��ڑ�v[�.q��3΍�x���.d-�W�'}�O�ۄ2�б�NN�A�w�.	�?;�Ѩٞ��-q�F�x�h�_��t%=I?��IE�}7>���>_ۘ#�H�!1,\�K]���� ��}�(��1�Z�:�
��P�E�h�̰���ض��m2-Y����z��P����-&ݼE��I��̺�,nF�8���77�^H,�/�~r�2��Dqͯ��-������ra䷁��ǧ�:¶uӄ�^���00�Y�"l�cY:Au~��!�%�­�G��ёh��lKE�ą�:��y�H�W]��1��
�e�}��b�~˵�$(�E�y�f���O���Qi�+%B��>��A[��:�RM*�tnd�n�m�of'�O�6��"|͔0�ާ[�8�������م��(��@M�lF��aW���(0;ko�r��-�>BD̡ S81RJC�=�3�#�7{r�rM��^��đS0��N��炬��$�)� I4ؾ�ױg>!b�Ķ���IDTz�P��8­��6���e�CnS�g,�_���Z�S#��'�$Z1>��o���ǒ4!��@�ApאV�<P?����y"a�R���F�=�GH�)����� 	Rv�6���]����׍���w��gZo��^��g�x��}����G��nU8F!�� Q(8ׇєzwV�J1RL�����Tl�_���4D�om�u�)zz��=����$���B�w�˿0W�o��(��@�Q>[y%��:i�[T���E�8=�3�%4�5H�< =�j����zTP�h���yq�c�G����w�O	��1���p����!G��Ƨ:��B�Y=ǆ���������@Ӡ=��ʨ�
5�D�=i�*��"��1�'7���Ϫ���8�K�A�6�R� =�^�Z����q"����zx�p�%�*C�	B?�
��v~�T&4J�)��4Qy�镄EA ���cƂ�	fp��wL�T���� ^s��2M�Z�*I�jg��/�.H���v�qo9~8���Dɜ��Z�sz@g���-~���_���(�J���߬b%Ԩ����=b@s�Y�6�|@�KB�I��]O���������>,;��֤q� ?_�p��s�~��E�t��r���p�� ��^�������e�Ƿ�`���s��kZ��g�:R�[t�KP+��#��fm!��~��I.��}	UqW�w���5�����3�p���u��-��G�_�&Ʌ���ftZ�=j�{�Z_\��yy�V�eE�!TDE� �c!߱��MY����m~$ME�����Հdz^&�?|[ ��Yp8�5,[���@@MUv�Sɝ��`6��C��C�A�]va}{q/�pрB,�Q���-���z�����m�i4W";N�f�͇s=Q��)0r��g�yp}9�W��dL%���u�}�����Y���cbĝ4�?��P@��I	Sa�'�妢nE��^�����]���W��m��ڈ����*��R�G|��"G�ňw�N�m"1iԾ3tm�\w�H��0�Wq�r�,A\�C���sY~B�%�&��'u��S��r��79>�2��F7n����Z�>�k/�{�|��`�;^�p�֏�T�5%闪Wџ��*�F5�V֫��<���r��-s˚3[�DͻM�Ɂ��9Y4j�y�1��>ϰ���b��L��P�)[6�	�2�K$]�E:��Fɇ�s���gą=.p&0n�C8N�$���I�A%pѵ�Eߌ�����pڏ4l���;X��MH؇s0��)�
7+��u���.�̗E�S7w�%�-���E� ��E���Hxfҫ�yy]��̚�R��Ƀ�f�!�Qe`���%�q��[h쎚>
����z`�<j��1�#R~F��W�� �ΐ3G}�ĝ�A�aε�k�!a��T5�5p��~�F~�^�g�g's%�1���N��s�LJ=���e���޲}�ٰ鰀:��a�?�gd��z�� ��y��y�E��0W�D�Ƕ�HA���o''�u��[�*#��}1;�=��Fi5V��0�K�D�^��%(�	iF�DzZHϼ���&!����%&��RT+��5��o�r�=#},]�F��b3���XS�Apê�cM�q֢�@כ}�I ���F��B=h[�{ SF#?�ވ:`�=��.	�-&7dm���ъx=5L!��J{��!v�{f,[ڎ��9�@pJ�_�o��O�@xc%���Ɇ@�0A1iZ�k!a��}��!�;�0Zoy̅�,J�t�>���#<�6��o@)(��k���֋jQ�>� �3-�x�QUakJ@M#�K�eD_�#r�=�0���L�,�oLHú�1+�<����<�q��Ж�H7P��x�[�<,���\���hix|r�r�d�\V�ic*	�VI)�;;��鹭����	�>���(G�Mȥ�cP�W�\�CÉ���,;B^���]S�|�>��5,:&z�Z�+X
3���r�s�jsO���W�x�}�Ӻ���f�׺1h���p�x�U/��!ė;��(Q6W]Y��Xm��-�c/T.��4p(eG?����B���g�l�
R��[�&lbڠpr�ː���ջ��C��`���2~���`Ác��W�d�X�p���QƌW��u�[*w0-z^Y��-�dR{������ЏAhl�e]�cq.Z�rN�����
Q�rSݪ��/�UTk�haq?O��۱��ӿ���)����!����(# ��� ��:a+�]���f��wcm\�m��N��Ц�İ3��ȓo��?ȵ���((�~Q�[_3�&�uPŘǺ/��ɾm�r�L�W�{<�>JQ��G��A�_�f0 ItxĊ��w"�.�cw�
U/�����h|� 
��/, ��U���a������D�`���T�_ટ��������,{x��z����\0%:�[2��ۉ�?�衟��Ѩ�[\Ì?����4P���<&���s�k�pj�AO���l�J����m�~������(thv�lL�?Od���\��s,����c��Ϯ8� �����`�1�N���k�s�Q(�(�BR���y|��2OP�c_�<��j�`K�<�_�a�A_�Ă3���.��7N�j�ugT9���X���h�]�udN~��ɀ��������`��9ԴFش��k#<;���	�� �u0������f�O�6C���V)鼥��X��Y:5�cr�ƾ����s�� ;0A[����T���u~c�,rڕ���T���@�ƺ@��)�ƒ,���Ԩ*����&}���|n
s�X|�G0+��$�x��t�{��G��gԿ�T���_}��3���� 5��6�]�j�a�sE<�H�i�����͐�q'7B�=3ƞ�ff�僐W2�s���� �[����;.V�~��Xq��_G!��{<r��Nh���䦰/ ���b7`��~�m��Rd��gs]�;�儸2���nj��$�Lu��ݾk.��!��4���C_>��)�F����F}�`�7��{m�z�E�j��Ӹ��u��cH9]l�b[����Vh�,��lFIv��ռ�N!mm�c���#�G���=�~�6��mk}�`$�p�D�;i�>�Z5�����:�/Mefu��Y}���}��'h�7���1��e�)4�I$V3ve%�����x�t�-� �����U���$���vڱ����/횦
�����o��0mi;�Oy�Vq�f��iɒBZ��̆6��'O����n=dA�Z X:�~����ߨ���/�	&��7sn%7�[6m��v^��]5�E1x$�2C�DSg6�d�B���iP��JUb�q-/����O7ٙ!���	w~N,+��5B$β��zo8�'��6�|�,  ��m�2�4YY���ht8�cZ���~Н%.#-%,"����g˺�"J�׊P��^ �ƻ *(u�(ؗ_l�Ծ}�J��*�?��&%;#	�.�'�G>, v� 5��f�4:�(�b���h/`i��� ��yT��)Z�Yz��=� �Lx��(��*[?��'�����~`X��`���at=�f7�7��~�k���Ow�5��U��c:,@] xOR�����d������W�:�$Y��ߗ1r��5mn���%�X`-����;�{�C���&j��ߦ�WH�s@��t���ז���ʩ�ѡ���k�"$�=9M?-�K���9� >�"�s�����	�����"�h�zKS ���$������j�ʲH���1ϊ���;�-�50me����Wp��ą)�'�ф�b���a���}�U�ENE��
��(=��P��@a����Ҵ���h�;��!5Ļ2�s;���0R]R�o3���e��܉��k/�3{/ZQ��Zx���_��	tV7�-���d$������Un��J`����?�0Bw�o����������B3��V�r�l)Rl�T�zt���mo3$Bbe��C�����"��:����ʿ�p���I�r��7G`g��MU�����Gooϱ��𛾦%�K������8;�:��V�/��?K�ntx)�3�~逾�GApB��dT�Q����v�.\�aQ�@TuS���&�X~B{M�60��R^��	߄��-��c����(t��Q��[���� t����OI�6�p��YPۨ�J�Y���5�<];�Y�
��H��o��\��{@�����>p܉7ts/�=�S,+C�� weG R-�!�.Iq6�G�bc�S��ŖE��j������ܐ��쟧B ]�U�𼱽0�7�n������p�3�	=��e�s�%��J̸�Φ��a��K�qZǷ��W>������E��D�e$:qVz�+�z��A�zx@"��]�Dm�CРm���/E��*�5���k�B���v��K�� o��C(���a�;���Y�����f�G�۳�������Ʉ��=���}j�vy��O<P�5Az��HG}P2)�yT���oI����>8W��h���s{2�e��T�&n��T��P��ȰI�:�V/_�\'���^o�t ���=�*�jH��.���O��D���l�yv��O���)�;'�IGeEc�U*Q�!/X�ᵤ�����P3�2�\H3� y���ʓu��L�?�R�`�x���,9#c}R��ڮ�eݬ�b�b�!�P���
���`�
�r��G�6z6� �CE�@= ��pT�� �`V�_L'���{S�8OŬv��P��,���n"�)�Psb`�1/,9(˲�pFꒋ�G�q�M%��M�\��0���B*~jZ+�N�4�i_�9��fQ0�S+� ��Ρ��~��V:wr�����*�${�w	! �������V�&��}Kڇ�i��2��S� >̛���%������UD�vj�⚥�okN�;�8ΐy5b0���1[���m�����.L�vq79�/���Ypv������#�������V�u�sy��1�!E��j��xe	�P�h�0��6$��+[>b��p;18	`��xXI��dm��570 u�G-�Ĭ�P�G����(>Q=����GPu��*�R����D��[6a�X�/�7�����7�if��0�A
����>�w�Ω�o��x��n�����D�2y��٨�q��J�N;���!	+�B�i�û�$�a�W8tb�Q�t�[��9��'����Ixo�a&�n�CA��j\a��4�PsŽD5bz��G��f�v��t[O
�ָ #EH�=��_$Ā�&�	����|gķw��j]�&ȿ�v'�Iw���S��,�M�V/������H��pB�p)M��[�9_�n����51�Z�T0pi4yZ*���%����W������Y'�K.��q(|&�S,3��b�����������<��1/h	�w�VL��҂�u�jT�pQ�b^���;h)��4���7)��z���Io˶C���K�Bt�11��I����rzINZ��aM���)~��WG��B4�������Ot�MܤOƶP�cM�/�����E�| TzeSu��Dwlq+�16�r���GW��L����tsupP�f���$5� ��98(�����������!^֊"�DZ�_��1���vK�-t=�9f
0؛�a�QT	��V�z�m�w�0���wbV�k�%h�󡹤�,k�B�v�����;�D��v�d���2�G
��n��Æ���*�ӱD��(Q�wa.N_8R6GL8�%y�hsB<^�T_��/�!�d���=�ϨM��h�h����$�~�}���]G(y����NYy�<�G����/�kC�F�قD�@>�ظ�������}�R�myv���6v\(�^��>��[1�wQ:���'!#I�9F@���no��y1&�F:`<��k�y��n{o����ccd���G乢��?�����]o��S�o�K!z�L����gg�H�L��(����&'��me�d*1޺q��N���Z;�R��$S"Y?��p!L�ߪtyx��Ձ ���G�Kpj��Q��נIz�0�Ep��*g����5��^�Q�O�iO{�n!�u�~��^�!�h
��?�R����T��Df���ñZ"R��S���5j7�ws�LI����Hj
��o����_��*��v̰[@��	7T�\��jf���v��֛�g�L�.Z�	@8�m�+��e����:�r���b�f�P,ŵG�]A��;�VyM�\IԷ��}m�#��m3:!�S��ޕ�w7")/U=��-��xӞ-����u����ݿ����2����HE;{b0�Zl̷����~㛜�+���!DCx	�h�ǋ*ݞ9��[�1�8ī�9O�������ƿt.s��\�Ѿ<��x�g�LoY�іB��<��©7��'���_�B �J|v�I��rG���9�"^JW�i��Z;���S�B�7�bP�*yT�ae���>-�0֏��W�G��B��g.Ђ�<�L9u	�~G8�	����-�,���g�0�}�ܺ���UWg��Q��b��)>��9�� -�C��Ҹ�;Ɯ�5b��rvJ��@�Q6��EEW��/3S�_0@���21h>�����_S��#�I��B�����
���$�0��(p��qztT�?!����Ko伜s���������wy����ˤ���iZ�`���f���ψ��<�Y=K����c�y��H���k�g+�BU�]r�5�q���NT{7��o��}�v"��YS9M���S8�k��TaM`�y�M+��1mźщ���E,�"���O�W�%YKė|��}�{V���;�7ђ�.�K[#�3v>A �eT���orA�ހ5Q����q��6qO ~�u����;�=�:Y:c��jwۏ_���S(��-�y~ 	mNY��m�~Ecw)#��������eۅ<����Մ��s-p�y�Qac�-ftw�P;��n˨g�
dł����htW�4�ٟ�A6���	��Њ[�&�wk����:5�Dq偟��=��8���w�2*�K���v0n���:��j�
r�W��I	���o֙ #1��m�8�Oj�{������_C���rYEi�F�y�J����bj#<�^�.0Q��ޞ�y�C5������v@�1֙��Y-�J�2����K�\��3jV�MҤK�3ms����;FA��fҝ�U1(�.�+9xW,���{�@|�u�[��-��-#�s�U44��u%\�����d�f�a��cE��9�F�.���(�7�q>��=�N��̊��u'=R����m6�\��%1u3��[�]��θ_��!��o��Th�02-�.	�p��N0��Xu� �Z`��g�g��T8&��c܂+R��kd6�	����To�aj�$
xb��@`Xʞ�\��,/>���WX���w^ϡ�s�o(=�o��]��	q�r7�Nk:k E�� r[�i��./�OY��l|��$�~l�],d}�;����U����K���t�徭����d&�~���}���UOi��n%7dίn���>p��D���p_�����Y���d�'51��#�P������9�
���8�>X"��V .��� -�t�pu�o6J�s�b��|>_�-4�!J^K*��K�+�'|(x�b67d��5ڱ!�M����p�%�j4�J�ʲ���Z=�]��!A^~�Y�o�a�u+�c���`�?����h'������%Շi��Fvɇ�H<�c]uF�G��_fU�U;&�ɽY��Ep�
��Ȅ�����9Dre�ݟc����! ������R��_��z`J�B?�Uߔrq���b���%yρ�i�z�gb�.5���5��85����M�K�Uu��lG���>$��pi*cs�سM��@�,(6��5���� �qm !�"�_l|Yx�5��s�C� ~�q�|V��n���S����a���f]��
#��б.pTu�Y��,D?U�8,qg�0���I����'5�]g�n`F ����	�`f�B�h��F���8o�EuD��̃*�r��6+AUdz���BL�\�w9~G3���݂g3f�A��y{�v��lf7s���^�i�O~:Z�Dg8�-�͉?E#��cM�<uWࣳJ��Y��,�`>1����r����/�'g�w�6�ܻw���7g�m���1X-ef��Fx���'� �dq��j���f��8jl!�T� ��:1��<��|�0�+��$�%�H*8������(�YnH`��S�ֵ�c���D*�x���y1Ȓ�f�7"ʹ'�J�*x�,��M��&<.�IҐ�9i���������,�:��x }�mqqS��^�K� �����y����:���S��'y_�h���6��}e��d�>����(�����=I9Vk�������3ޕ��Z$_����-	���Wu�a\H4������E�?�z�Sf�*�%W+}��=�{����AF<
y,(��<���`´I#�%2*�[She�u�,���C��`C����͋)d�5���g�v'���<A�0&ߝ��qB�Zy��� ������NC�]�0	9��*�}�|O#�%���AV��Gx�
4�9����G��o,6r�W"��[̸�!@費2��8C�:Rސ��p n��並{��b�g���(a���Jat����F����:Q�5��L�˙�2���ˁ�F���B�!�u�8�#w�͜� ٚ��nfs>T$�\���^�*�x�G�����a^������wѻ�Y�݇�O\�̅?�)������sP:y�A��`�W.7�0�����U��hW�Wᗟ�Ŧ���Y��̹U�>�~��e �{=�� Q��A9��"��SM��-��Y��=)���[�5����r��N|�NAu~�R�'�&�yK$�lͽ^���I�~�)��_f���f-���C�R4d�$�1������:J*f0��>z@ �*��y�jz�nG���#�7�e�?��r��7�FGѠiW(U't&܏z5�jVu "^��7�]Fܻ��#����+�Wn�PJβ��ƭ�e�c���{˻Կ�3��=we{�tCD`�����'�5�Q���׉�O��vK�ob{;�Q��_^ZtY�o�'�r8I�$���2�_�� <�?i̓�I���-&h�'^Q9�C� ��>Enwub��Q��f;���ҙ=��*C�y��u� OZ���H$�GKO��; #B���GA�P-$�q2�T�V�QwD8i���Ni0���#xT�i�����"��;^��aJkH�sZ�[�\���*��y����A{�ϒIL��T�5 �2/(v�d2SD�����Sp
�/`A�3�P"��jΖ��,?�R�oWG�'"$G]�{�j;sH����)����p,,���y\X��PEr�hXM��Q����dN7��
`! %����b{��c�{yu���=��R�$�OmXUh�O��rH��������.�ū�Ĉ��Șxq�3WmКL���o}��Q�a�f1�4?�S�EFm`[lAs� ��l2S�y��J�#���yO<h�]1�$,�+>‪��͆+7(�ʩ ��s"5�Ye'�i�P����iC4l�޶ўVM������3K�"����!�?����~��/�섏��9��&[��]T��򇜾�Ӹ�x&B��MD�+�ԄC��S�n-�f��T��O0�0kE�B�*�"/�_��`�}�vժV��U?��C�����6x����m������C��Z�N�_��G:��c$(q�Q.���<Dw|JH�H�G�L��6�a��0�t�mQ;񏐬9�\�ᰦk:�R��qm��3�R���ډ��{�|��z%�+�1�1Z_�� `���[��%�m����L��"�?�J�wd�C�2�b�2$^|#c��d	�jݭ���UH
��Kְ�W����������I4p���	���P+r��h� �2ax�ԇ���'9m��GtRuF���0F|� �r7�nQ��)n��$�$WS�e�%J_��n�L��%�fmO�O���2ȹB�J�����1�ې	�ޓ�GN�&U�Ճ)����aV��Vv�� �foj��Q^�ݒ�q�W]��TԊ����H9m#�l������?�(�;%�f�F�U.8=5{^𝵭����K���)�?ʧA�[(d�*�R��ٞA��T͐Oz��@L*��#���8�&o�+x�f�Dq�rЇէ�upn��.�
��ך�Fn<VU/"H8�l�:B�o�V���4)@T�{�!����z*ͪ��?� @�ho�5"L���T3Q7W�����&���O�!�8��b{Sy]A�h�`��K���s̃��~$.���|�I�	y7rj�xcd/�|Q�E'0%k���&���w�0�_+���$�Kk3L��Õ�w*U�d!����A��!I@��髖p�B�1�/_��'����zQw?F	�֗�ݠ��_�xfD��1y[���"�-b����乸��${�HY?�]O]��~ۋ�����-�ez�����
����/��IcRM�'�K4M���v ����h�l�Ut���2�||e��9�[Ne�����(�9y��!��(�uI H5���� �7֚`�u�0#j-Ű �p�ch[�IRV7�#�I �!����.t�i�ߏ��sn��$�.׶�R��c	O/׽>h�(���D�5��� '
j��A����5\�R8����j��1��]l�����[��R$��] i6T'&t���R��9S�Tu�x+=+�\��1I1�J.���/��%:�����h��?�/p�A�v�F��Siӱ���}q8eR��
F~��ǎ�.�g	TĎEO,2}��x]�y��PΘ,�K�8����N�َr�t �&Z��������r��__o�ב�
�u��J9,v
�K�̏����,����]pf�yA��Pb�AF�M�8��%�9Z�0#���o�$$�Xx ���S���\3'���M�V���@�����0eiMsp�-���"#�� O.����st�v���.���"w��j�)�.k8U`�D ���I��ؒ�Tw�(��g��5)�Oa�=�̸P��%�G`�����B��W�M/��Y���NIuD�	C��|�ϸ/�c���"p_oq�iF_Q�~�J�Q6L�]�֭6zϨZ��$zz�pT��!	����ԕ&�|�;e��1^��A.����vSf���J�*~��#���:kz�U\Qe��P��Z`���!��� o��b<���%��W�C嶯�\���,�ԇ��C�J�i駻��@_�) G�%@FPr� ������/K�p��G�p�/'��Er�ݺ�|�5*� +�N����7���Hsd���?��֣(��ɝT <�kx��xhq���6e�i��v�7������3��>�>�uC�Z"��b�����0N}9�}(�}�s4�RP�.�rak��Q˔h��Mò-�/;��4H�,����O6�����fGx���MGe�29r��{O%�3L���F��@!$'+�8haG�K�dl��ratS;���bH�P���Zż��6zڐ�J�׭\>�ʳ�汸3���	��r�-C��$�wyM9��3%X�;<(դ��1w��}�#O���w���A����	�gBz�SY�rZO����2-���~nɧ!��D�eRu�ǽ�Tu�D��E@�V��&j��h׃���&�ֶyȼj1�(7��l����^�|U�9b�<L�����3<{��e�����"MV	�1@4�y�����&샱�Y<��J���%GƠ}֯R��Ď���Q�Y��@R�_T�I��F��IB��E�$�c�ha�T[lk�dr��R�P����^��1},J���U⒉�����~���ӵ9��.H�Ɣz�y�j���x_�w�d�mF��y�J?�|q�e��J7-���F�5���RY�.T�R���S�3ߜ5̮�X����@.�)
��q*�Q�.��qmp��UԲ�QWmx/9��wM������ZF�ҜT���Y�W��/˒72�#�������=�*�M�0o�!V�HR������x6R}���<��<d���S�cF^O^"z����%�o.lG*-�#-�NyD^�!z�nM�MZ��{��׌I�i��r(Ŝپإ�s��YE0�be�0I-���"��ي�Y@��:���i]�O4Tլ��H������}i;4�\�Yԝ��T��H��&��g����%p2��$W���@dQ�9�L�[7p�tي��,gpf��{����L�!����dD���LN��]=�s�t��.��;)됒m%��.U-���Y�|8z��W�@�d����d��av�et,���u�X�.��v�A���c�ب�� >�$���`-lt$O�FCNɉ!a�쭖�>$mL�k�yr�c����:�����-�v��]�T�"6)�r�~v'�H'�Q&�
�����GM%Ǆ��$�Y6D|��*�q/i�It����<���ih���8K�Ԅ�R��>��')��΄Î`I�m�T�[n����R�,�,T�pb�wlK�˕�4�c�Ց/{\��T_�$P�x-��'�;^�ß��}�Z&0�*���.�^� �������Vg���f� ,+�?��*U�����31��hg����ΰ�=�l��RwS�F�M��S0�K���g#�짋X��'�[�E*���pSx)g�P^���M���F��>���xw�㺚����!����[f�7������O\��g�I�p�67�n�H�oE�׼�H|Z�k
���R�I���u6��]�#[ӄ_��9�ַ�S�bꦗ�����^�0�����W�D���5�(���ΗP����F�N���VN�
9���#s���h���F���4&&������ܥa�cv���!4aOVh]�lZY��@Y7���**�G(h��`d���;�.��̾5��6��Ny@�ѷl2�voi>�fz[�Q�������J�t/c�TFن�S�E������4��
9�t�g�N�"G��k=WI`(̙��7Y�x$��.*g���D����1GN������x$>㺕�\��<�_�.��He�E݉b���;��9���Z��'m��,:����n����KE�W1&bn���V�t� �ww]]���9�P5YnN���{�~DT�����
��Z#^������EW
�x�uA��	�}�����E`I�3F(PCFE޴���P��x8}���d��ۙ��Ȟx�7"8PN0�4Lt����b��L�`č������P^m�L�>}J߀ت��.P��m$��57Z�=b��-MO#�80�V�Q�Y$!i_�W�������Js��4ׅ�/0s`��+���e5Wu�6��BMap()���d��-{�-�*	����&Q���b�s�m����16���I�y�E(�2�Uz���-�#y��C�YI��PS/�,�H�;a�4��
1�JcsӠ�ks�������@�.�:WG/l9����*���\/�O+I�(ˏ\M��o�(#�!�^�_�u9n��  =T.4��a5�K���Oq��yQ��^mr#��ՓM��tW�5��s�Y�N�)
�r�߹L��� ^�a��_BL�+�Q5z�_��
ۧT� ��7�O~�����*��v��0�+�4zc�/���!�v��ϕe(Sq���w���!��=�.� ����m�z�q�H�W��8nֺ������˕� �#xv�|&�������_\�M4J��X��/�h�x��%�+��9��@Nrb���p��4b�x�|J�\��*r�m�xc,5�"\Ä&S�x�TQ���#�B�eKK����Ӻ�
,��|z-����;&Ay��R�7�a[�ˁ29�������(�9�-R��)�ug1cCy�n��Оy���}�1�5����Z���ϯ�\m�N��E�Y�
o�Y���|��]���`�9�c�=�)�0c�I͐�Y�5N���X�l�+E�����)d$D��o�ؓ�����z�-G��1/��n��~+.Ok<�T�B ��O{��>j�F�I�u�_����5Hl�E�<g0tt�������?�tx(C�+)-��a x�.uz��K���
���t1��ý��@R�g��N�x/�=a�u�#/��Z���̱��K�~�/�Һ��<�On�y��ZH�=�}��x�gK$��OU �o�,�(=}O�T�Ph�\5����g{��G��L��B���`�N��ٴKr�9�jv�@�2M̲{���Y�.oó�h�w�=}u��$#F_2s�\�C� 4�F	@|���]�_ݲS�`�	7����r�+��TĮ�|����jh���}����6���z�m?��%b�����zzGy=��[;�3����૿��C��������� k�`�KP�C��&� �����W:/Ј8h��C�+`BQ��X�rԈM� ����F����jU3�R�BX� ���8�6w�7��լ�D{�(?�w��.�<X�i;�e�`��z�����`7ۀkmoN�]�[��&�$�H�wӟ>�B��]\������yX�e��k܉b� M]�{��J/	9]po���_��)��v"���]�2R��T\^I94w3H	��{Ul4\����ݵvLtw��[��:���>����Q���o�n����I=�D=�!}M�3=);��p��c߫TҾ�NZS4'������G��dk��U5x$#�_�"��6�Hiږ7�OC��g/N�<N�dQ|x�B�O�ÎZ9��ƙBH��E\MG���ȵ{�Z�.�[�pV��#-ʫ�W]�z[>-8����/����$�uXޢ!��Hh�xٵ�f�,?��)of�(&�J'��&�X�쇀��A����� ���=���|<�v�)D���B�1|��*�;���{{�|s�i���༈��HᅕĈ�z�X ����Ֆ�4�-/������kk�:�Z/)��m�<,κ��oa4�բ�98��Fy�7�T��/� ����Eo��%;�oq�-�7c�UL	��ҽ��J���R��?�C4�52�K�L�1ϳ�@�����|1�[	�)��I�!��������_��s/ˏZ��
�F�4�	�	Y���)���A�m-��u�T7���2�
?Z�>������"S�`�j�L�'��	a癇!8L�g��8�i��0g�<�w}J��R�Ww9DP4r��4OZ�"���ŧM����{7v���W<�O�vh�ɤ�Z���i����h����U��Gʆ����^��x�����_p�K�tL4�ƥ.�_%RO@w���e%���b
#�Ն({�;(*����2DB�$�/���s���m�aCk�����I�g�B�4ji�ψ-�7�v�?�Y]�C�8_G��{#&M��91'�?�+yq�XU��Ze�E(-#9A�)�]_~��[v5郼׫���}]�X��u:��
����I�*�-��_�h��{Do#�؇fw%��E��X�μ��A/�8�/�D���j�"�� �Ž��[j�
��f��X�z
�(*�:��X�cJ p���Ve���	5���#����r3����C)��FZ�źOo�Մ]�T���@�{�u�4l���˲ �c$�7�^�3t�b�)�,���1aL�����XÄ~�ך��F�v�2A��]���uK*�(���}m&[M����ِٜ'��(���w��A�Q�|2Dظ�u���p����a)H����0*3A�����~EZē����=�ŀ�*H�[>��+(s�(	:l^� �h�<�æt���.��cW���g$�?�H�2G��E[R19�!��R$p]'I��]�1�����3���9��������@�p������_�=�I2XJ���U �
�ȰP6�9�4��> �L��8.�3���^R�0g�ηqg�����[������Z�m�	F��UL&���Ro��Tl[;00$?)�������8�l�.Y�@[W�b���P�s���*D3�i�X�<��g�>�O�CG9H�n]��B�Eאh�7Gŗe3EvG�1�b����_J�����{V'���G�$Dָ�r�}$"F�Lxd�p0rO�������ά����x����8��ʾ���󟕧-��l���E�۝��<�װ�5 Ym����_�U�Q����|5��O�ƃ�����+��� $��>��m&̉ꈧ�;��[��p�;�$���Z��QQ1SM"�ش��
6
��!vެ!�Q� g璚<zXcRP|��̠��4I~��я�W~�8r2� ���>�XM_y�!b�f0�S���p  Yy�&o�>1[�%�V�UL����q��;S̺�+6�SI�}�0�Wf����O���[}mC2���������Km��L!��9��e���7��~l�{9��G;�J�����&dM��HJ�5��47/� ���@e�$���#�"_f�_&���(�:q+�7��&"~:k枹��W4�}@9����S���|�A���
+� ���Q2�R=�>�Te��t�����>YDo���s6v74[�F�x�'�T���^�g�PvDwg�aSY�O���t����>��$�`��'v3��fs�T#�OHo��*��h�Co�
�����LD7��Ҹg�y�h	�s(E��MtE=J�i�9�J0B%|�|YY�I�	���|�����4����L�7?x=�<��-�"Νc��f�~�i8O�b�q*}��7N�
� 2�'�o�P!5�l��,�H����T�估̮B6�#T6�������:�$]�E�p�`�4 �E�Ն:���\�dY&�{>�������0H�� �x�3܇�;�W��?���lL�����T���w�"�����]m*��kR�V�Y܉<z��m�'g�հp�����C��l{��p`���t��|����I���������`�q�(�
%v��/���!0�3U�G�(�g�� u����&�sdV6?8ٰ�8�s���n*�U�@j6FO���pzQh�L�!�F�p���To�tz+�5��ԇ���6�	�M��	(�Ű��+Э�s*X�ц��`�4���3j�Y8E�4](F�7��������g���2Btﴷ7y��b����ZmdVd�2�`�îYG��5`*o�ư�3�*	bgX��]=�3�H��j�9�l��a)���x3(+ 2V� �+��=>���o�`�w���3�-~��d+�R��ѠU-s���y�q)ß���TbX����mbV��֡g6�.N��d�X]Y�N�����N�h9�Ҕc��`�W��P(�e��J�:��^����t7�.�<T��ݲ�<��P�sp 廙��xS8!0E_˩1�eU@Ә��m�Z4֪�"�ۘ}2�I��I����am�V<m9��=Pn�
��bz�Q�81y)�'��� �F��#����)�JF�o �
(��,�\,T�i.��Z�v=�\]<���j�s��
/|}�.����:������<9����\wt\{���#R���㿦���K�{3�|uw��H���R��w����=�>�%Ә^����J�Ù:��iH5�2��1����7"*Ջ���ehRcElL���H ���t��
��5A��O��l|`H��"�h��x/||P}٠��6���k�N@�T)�Y�h��)^�9��q	��S���CS��p̤�r��2�K;/�)i�O��<��ʵ8�n��a��@hp�á�W;�H�������/Z�N���}��O���=�����ۉ �l�aË
���]���G������*�d[�wZ��8�k8"�m=hk���0C��5nW]v��.�'��gj��;�qI	2�EҶp��A#�W.S�9f�bA��,�07¤����m��g��H��2:�uaCtܹ��V�qb�{���ے���ً��O2#1�����<�T���m:��v"��y�d;�}fNu1��E�QK�P��7�ţ��L��~Ug�Ɛ%&�⯆/|��ޢ��ˏ���v�3e����#�4<�xXȮ`�k�4��bpm����R..<+�]E��z0v�pSDb�Z�g�Q`!�ioKB�e�n"U��|BnMURH�B��Z���m����#fR�������yԘ8"����@��g(+�Q��{C2�Τ��Z9�*�ȥ��"X&h��9=����>�G�Ѫ�9}�DD��l��#�L�}���NP��K(v��\{��S&���~O�|%���c��lr�MN��[�
"D��{\H�<�L4�o[�.�9;m#D��-��EŘ�q	%���D-�Ե�J��+�+%��XY�]y��f�� �$l@u��]>�C��l����J���)�S ��Y-�k���ҏ��?���S�ќ<�`
�7s�_.RA{oQ��e&R��?���
���a�괻�b\����=\�K�5{L3��A��0ў�3\P���'j^��<#I�L�Eq�;T^/���.aw$��6鞡��T�k�	I�pЏ�0�0���~Ȕ�1�uޘr�'7�R���~P��ʅ�m�N��^�9��O�����f���Hsb�I�#�M
��}r}�ќFF�N	-h�e��۱��'��pa�i�R�Ӥؒ3�w����!C?֧tAPҀP����B�;4�!��B���>��Ȍk]ܭ`b|�#�J6n���2 �<��s6�Ӭ@�Ɔ�oK�Tr�-g���?+���<m����60Re���r����� �`	�u�A�v�8^�ެ�UZ?�Z�� Qo&3������Ū��s�i�W�0u��X��)�E�}��^���m��ZE�R��y�>�#<d�R��m��Q������)73��t`�h��3�GL�x���Gd�B�o�Q��]A� ��kk]�t��J��Qg]P\8�������{��D��̴�Q-���(.B49V�`�ji*nǿh���6��z�q1��߸����<Z��_�ha��p�)g���<�U�&��Q��OC�#e
����t�wZ�Nb��T�?
���~<�C &� ��~�:�����b
�2[�~�����Ҍmu'@�](p��8?/�N�դqLeīAHD�l�:n�?)`��¼�Ƕ ��y��;'����:w)���V���B���0&�����U�����$����'��kLt����;��I�AU���Tͱ ��W4�Qy��f��������׾}ˏ����������L�/t�?��ia�Y�Ȁ����Z3=�p�I�"{3��:���`�WNc�%���o���3�x��"(��+����=T��I��,����0qv�R�Bf[V�?���+����A��xJ�N)Ht�I��q�ۑ�V�P8v��+-;�}�Ą��c�3B�E$�ĭO���c���!�.X���Я�s�m�ć/i���1�cL6Rj^��-��G[ͯ>���NM �%��������1Ż��M;��^��V���2{:��������@b狀Ji��<w���tm�u�����9x�WܜԾ���M#%���}#~%]�_��wS���Ue
��-���A�:l=%��{m"̴�R)x���t�w�U˶����8���;���WEj>1:�gO�Hz��Ml6rn%!w�0$Fp���p 
Kt�rt7�h��q��b줇ō�`b��Iz�Q`�f츤3��m��� �l��f�|KNt���!%[j��r`������G�޳-��
��&0��'m���Z�[�Yk��ѳ	#I%p	%��H�)�c�نk �zQΌtX��'p����a���j����w}e�����ɵIx@HϿ�-�w*ph�K1�wV^cX� ���8�?�ӕ�A\���ty��O*cŤ�l��}�����63�]BC���0�ǹ�
���;NX2C�i��a�s1����d�A��0x�_�+߮?jͿ �O�>,^T��ʾ;B�������ZU��VK�y���x�n�m$�0���t�p��sz���1j�1�����=d�p��v�_�gR0�լ!�$%4�� ��r�����L��r��H��i��!¿�k��e!�n`ve�6�oi��!��(�x]�|FS�p~�@�R���BZ@γ�~���� �/����Mo��ɴA�Y}墄K���mMQ��\�+�%�u�|���L���!A$Kۦ��!}f��cq^_�kg�7��!Do�l�#�� ��p^�l�����B=\�1׺��?���4��s_�[I���ũ�X�r�A��+8m�c�����?.n���?�0o� c�h��l�.����#��K���ñ�O���q��F;�����yf6�TWl�m\�6�4��������[�_��v�La���~o�Q�!}4f�P٢����o�pk�V�CL'�_O�S`a��Du�)�3yĂtΧ��p����*zby�"���!��6�/E��o_�J[
컮���>�3L=T�ųa������-�.tHG^��'�����bN�@��m1�w���H���'���DE:��"�f��P$}5F5�P�qv���Q��yY��5�Y��Xp`]���4X�ޖ^W�R7���i�Z�fR<+��� s�?�Q�Tf�̙s�82Z�qvW+n�g�����';�nu=@E
��2sˑ�o�@=7���8�j�$�v"��P�w[����1c�W(�.����]���;�g�E�tB��!!-GX�\�V���2`D^��tNƴ��T�9���ν��5���oǭ���9p`�� ��_�d�uj�R���I��Tp���k]�4OQt3(fZ��q�Yp*�Oѵ����J�������d	�-N���������߿�{�<�����:5h���,d'u��.C��&F_��3ʺ���jX�nk8l�̓y�Nr��m��X�g�����Z�������\%�r��4�B(*<��g���ڔ����+��W�a;�
�����̕�n�5�[��j"`O��F��DA EN�0Hz����p�ty��1��]+���j�~i�����L͊Fl[D낇���_��u=Y���Q�:�`� Q���Ed=�e��k���R$�\q�q�n�PUUmjZ�e e�#\�|�ّ�Vt!��o��H.S�h�A�����K�e.Uk`���=�؋7�w{�;�i�6�S}����k��IT	��$0���fB*惹S|#�_(%bfzu�f�0�$�y��/9qHp��g_q�'�u;tp�\1+"�B��������S�H_����
*��R9�}�0ʞk؋�����.��-9�ē z�O��~�Zr��w@Z۝��ű����u;�{�J����%��k0@�d?���{G-qN��3Z��DW}Q)w�{���s�Kzl��,�-���>��T�g�u��d7�˦��OxP�u�-�gK^ڹII����(��x���Mp1йH�2�h�L�! ��`��F���ً���Ք8?����U�U���H�t�K-jsK'y��<\�㆟�a���6����(A�~�'D>��j�f�,Rk�۪���P�ܠ	.�2;Y�(S2hӽ���#R�ň��M�<������}#�-�L�W|h�5�u�W� [{:�&1�g�e�����+���@EA0�j��(.SG�n�Ê~׶�q�Ǩ.1mgw�t��R5�`Q"Q�Z�cF��d8�!�N�̬lv>Х�������S��̖�O��b.lE3���a�}����%Fhi����ެki���� n3��} '�	,�������$S�e_��%����� �4�;lk����7R�aF뤃�4%1��f����S̫c���MW@9;�u��j�rv�a:h������܆Ԣ��A�����s2*%v�
��/6������wi���W�
��"��c�RI�a�_Jo�
r�ERMe��fc�Y��5�<�I" ٹ���]�W�ߍ��"A�p�ݳ[��ZOk��g�&>G����!��9���#��n��(g��ء�4��vF^P��.���`6 e��� ,+�U��f��lɛ#�W|A ���[�|�_ٛ���XŨޮɽ�(�= ���^�5�14x���;�mp��B���L�*�$e��P(r���v�U�J�3u6k�n�w�}���@�k�[a�(�-뼐��nǂ�J.����_۝8���U�ګ�,_g��G�3n(����sG��2h+�t�޷=m�˺˒��JUkc_�u)����`#�����v^�@��@�!�3wx&�W�Y�6�D�YꚝX�S�|����D��m��9�bxZOn쎴���E�����8X��ox0i��v��o��O� L������\:�ir�����Շ ��� ����A�������;���m<C�|�����
����d�d2��z�f��ά́��D�D\��K;ڔa)	��[�l}�)�0v$��3Mk����sN��\Ԕ�E�]�I�=׏k�yP� ��g :�CW3�ɵ�����0�}��/,v/�]���*���l�>�}ηC���c�e��$R�c�o�ڔn������3I?w�x��YgN��ԈE͗��`�;ƨ�t���+I�
�f�n���%h����[Ou���T���(��d�΅zß4 �S�-�\�a����yU�t�������U[�&���hwu��iZ�.S&�at8�A)x��0�l�yN�a�+3�hǹp�8�D��4ff9�+}H�^�|�.ӌ�'X��4V���������"��������k��i@@bQ�g4��D���vz��ҐC�{���
��1Z�4��f:����Ǥ^���6�:�L�4C��J|~�g�߾%)X�������p2A�JpElz�*r^)�	��\��7M!�S�zM�4��݌l��-!m��?����&���i`�K]I��ftV�M�N�������6�\	C)����I�o����Kg�k�GYZV]�&�����T���w�V�0�+���9��:$td�M�'���@�J�ۇ����,�zڧ(�%���Q��Y��	�(j�3��[��t0r୑��kk��&�m�J	�3o�/�TQ'��@��iq������*<��X,i�����"���ڻ5��/��".�DR6�qB�� �_��ɉI�eQ6�/4�&�ه���f�n�r&07�BNRy���)�W��f��4E�E�$�u�l��LkL|D��S��Q�j�"�f1`UN$s����B�/� l�V����x���CL��K�[��ݺ}�XzIvʸP���6�M���Q��C����H��Rw2�p1V�,��� ���*��<�a��)� ����h%XUcx]��J�}sZyη��g�ξ�ZX(�W���Cs�����O���D���=��0pC��@��;�����ƃ�ob���F
�C#T�.�%KH}�<�Dky�"���M����7� �
��1��9ea�R�:mK�Md�W�Sّ�n7����T�uv��Q�-�!����ț�+zoI��y����(��*+�?�n'���U���L(��u���o��J7:+��L?a��ş�X���U/24:�j�\�Rs)�M��a�Ԇ��L~$�2�)��_3�Xk;����Q6�X�ke<v���f�O,'*Z:v�a�[��� ��n>���qbg��n�sF �e�c
1�VÃ�1�k��Be�Z�p�LRA��$�\�
����b@�;�<D�������W/f>2�ڢ����Н����"�W���b)\�y�����o|	CF,��7��l�n'�)�`� ����N�8+DS V�qU"�*�H%�8H6��� 1G/фA�:
�lZ)��AV
C�����/�˓c
� �'�}/���x�(MT�4��}P�U�c�=Iܳ���:G 5��g����{�f�[Rr�~6�f��G|�m:����� �+EK��p�V;�$�gJL)3�ݵ�D�m��3MuY��fP���I0t]�]7Q�t���4����%N/�S ��<2�tfC��䗟`ρqp�߄�z���G'�h�_݋�} �����ԟf4�X�9AZ1|oXl¯_ݻ[퍐i:���ɷ�Y��hʸ�Ψ�>�AѺ�e�F���`��s+_��Z����Y1=�� pV@�[}��*�ƯW�E!Lh �7�al<�>�0
{�g��w�q���_���G�]���UZE?Ϫ�o~��� ���N��A0[��P`QMwJ����b����� �[��0JR�D9��F������0Ki1��"1�g���9LИ�FQ�b<5$�>��Ami�߱���Nh.v��d�/��Y�{ y�@}+���l�����[�; �ϧ#2�QPu��ԩ��|)ElEr�b�Cg��R���xX�b�1�	�m?�QE������IM��H̑s� ���r?�
/��,�,cӠ��)^r��o�
��nC���Z��+ڬ7���������_��;|�{Yb�#v��M�f�����@��X�Θ��?η���ji�g@�"��U�q֪Y1��VW�1%]��m�d@ш�F^��D�R���܅�n�<�	7�����?^7�q>�'���#&�E��^P0U(�R�;D[H��pܟS�5s�J5�����jۨ�-I�<���Գ<?a>u ?-�T���b\B~�o�v����0�;$L2��yX�js�}�/�S@)l<��X�h4�Eܡ�QL緿"�p�|���1dN>ƿy7��/�]�>?;J0n���l�<	_r���b�8�6����N\|�*Z.�X��_�ԣ�;@�;��/�YJD���X�c��t�yƽ7�2�N�.΋;�im*��?M�#�4����
7�#w�8��3Ԋ1'e�d���$�Ӕ3�I���_�Vي[�+N,Ah�!Ӡ�˙�On X#whrXIԎ��>�)�Zd
� 9MXN-�8�=mS�����cΒ��(�'=m�)��|O�'�	y�#�}�a��3����XD�ǹ����QJ��J���=ʞys��x����D�F^wNB	�`��0L��s�A�g��_��Ke��!���H@����j�H����hq���������Ty܇����t��&�P���2!�w�̊)��`��=���	�^��T��W��:Ş�M1��O�()��F�g�g��+�	b:�v/m���4ٲX2wщ� �kN"���?g�h����{[��~�2�(�i��pe���{L�L��7pͼ�
��4��(�{�� ����B��aa�$Z�V��^:DV|��ܔ[�-7�{8��G��:�A� >�ɰhv�ū��s/�?v�4��,/�h�E��e�N_�v@����횯�>6v�T��IL�m0�Cde�� �pZ1 ,|��9+|/��{���@��"�Ihl@ F�a�(�k���{"{ݔ[�7��ď�z���˒��5,K��§�k��/�ƽ`PMa1��Uq �H��T��U�I�xPu?#n�Vm� ��j=�3��|����y�̓r�!O����s=�a��{+�v��|����%nEI�O1t��5l<��_�`Ǥ
]^.��=e& ��[�ҁM�۹��`
klR.�fD�-��W���y�;�����j��Rq$؁�!(G��Y_�k/�~�E!<O'HZ��c�N��|�:��V�j�N	����bj��QSu*Ző��<�M�t�zǨ�'0�w��Lw؋f)lҦ`.e��w�L�E�.��`����s�ߣx}���u#�2�z���#��ck�Nն�ѡB����N���%�ى�׹j�z+	F�z����U籼���Z�ў�W��5w�r:Y�{���5�)�a�z2�W=�r-�s.n�S�M�X�r�L���_w����O�x�J��2k�o?x-��f���;Sj"䫉P�V8���D�
l��km�17Lуp����ف����P�r�y�]*,�a�F�H����L٨@�U��x�����Ʒ�*5=.�;��	?,;j j�zˮZ���/�����;��jd
z����|���,�g�C�x�E�Z'�Ʒh)��#�N'���K*��VZqн�(��J����{g��Ѱ8��cz�TK�i��Dk}����U�8�zwk(��DؿsZ,E�2⯬"F"8:�ZW*re�$�p�|�5>�fpr`1в
ȳ6�� ]�3�oi�F�4��L�a���gy��%W<{��P}^��+#optxfT=�����\�sʥ5�\����[R�	�h?��W󁰨��|Dz���}'<M���>b����r�m�ˏ�z1=��n��>���G(�5�By@�ڕU�J�A���@KM=G[[�Wyw����P5+���0��)#j�'Ay�*]��ªm�R��+Iň�_�L��_�b$G�p����Z���L:�n�>�d��a͡q�%�rb�T@��s1�O�.T��[S#�
ޣk�H"��r��[��3}�+�����6�V1�����ۋ�n>ZABe�Ώ�a���cY(N;{/��EC2��oA~s�@9�����k٠�7��� �7�$M�W�#���Fм��Q�du4�x��lid��ޠ�ۯ
Za��L��,�2��ġBW�����!\+���wQAQaO2�~HԀ<�aL֨��o��N"W9�v6��Я�Bo^�Vs�[:�:w��6p_�sηaV�4����]��ëP�����#/��9Z�E�I����f�i,������
�vSF/$�s_h-�(���;�X~���"����_���1�Bp�.KB_7���A�����:�V]{�C]\��3�_\x�0�?��P��6����:�Z#c�Pe�ښ�r=��+ �a[�T�,H��c��/�a<���&���B�ϩZ�s��=I��q2+U��#�u.��t9�+�w���(A���:��0��o:���oI��lZF)yo���X
�ZQ���$?�d%�����[����fXٝ����Z���Ma��)V�K�\Nj^�~@�6�?���ȡ(��C�s�5��$nu�K%�w�Ǹ������6��a�$7m���w�t{jۗ?�J��.f�D�ge@ݤ�S�}�tS^�����炿H#Pղ�@�+>�	?u�s���E$�Q̸gZb'9$H��7ʧ��6G�D�D��@i�gOf�}�&��Or����Zy���$�J!�P�?l��_�	-�B̿/
���������{��2�If�Z
2�˨�j���A�T#+>)��g��}�+��z���g ۞���q�c�?ׂ<�5HdJ��jI�)w�J|+��X�s�`���k�_����yU~��O� m���ʕ(��x�(!��h����\��*q�~�T=c����w�b�n�s�o�X��T����_�f+�r�U��B0�`!�`k����ꍪy�إ�M���ʐ�)m�I!`S��	
?��غ�l����r�ޒT��m]�s�S���~j҂�::���T�q�H�����gc9����}rD��!D�~�
|h�)-І\: �l0CQD�W!���ɱ�
�C��]���iHm��� �r�+J蹈�7�r�c���k�+��<=.8ŕ��9Ux[����Ö���bp_X�Լ+�����Q�ƚ�lSb�WW\��`�P�]3��Y�wMPfPE���#���Z�©'�Qx���G룉8�x�;���V��z��[�&�+T�}�j����w���%+�<���j���MM��@(w����W�M�'״����!�q�N�5�7�]뗛t�
�AsG�<�LH��(n�I���A(���{༂�Zڋ��Y�1>ؐǱ�q��{��7�$��3�p��+�=UZz�h��(.��=�ƾO�0`��zz�m���O�'�S�徥�F�NC��[q�2y��h	T^���Ϲ��̏7<�ְ<�%SNA8!~~2����:��)�UV����`R�}iS�N���s�)���9.Ay���C{���;	:M��<��vWy�[�e�#���l�1b�[u���O��5ܞ�M��+J�,�K�H0��tc�(�f�ae.��)�d�J���ֲoF�FU�6��1h������0�2�XcF\�
��kC�\JAr�d���o�@�9k�
++��I��Ч3��A@|,j��"�\#����AޱH�^}>��#S��UN�T���4L�����,�J�`�-�XiN����8�wh<N��ܴ��e���o�d�jA�]��B�O6�U.e�o)<�a�*jF��������0t*�GY��(����N(�wY�0cω�<٠���r��clzp��cA���D�`��ӘI �.Y���ʕ~�p:�
�P�z��݊6���	�H$����ד�]�{�As�\C����i��W^�T~L,�7�*��QGR��	u?^��~��A����C���a������Vx��r��U�v��.#�� ��Ċ�_y��ߕ�$�h����)�)�+i?#��
F�ʪ�'d��ûLQ�LwȰ� �J��Wj�D����ÙKOx�i���H�@�+����̔?�{@U͙h�iz^�'���	��^��l�uO=Y��۞RaJd O�B�d�(�k�1�6Yc�Tᆜc�f;<�;gAކY�P�q
�c�&̊����Xԋ<͵x�n�*�'@��9�x4�ą%�nM����!`���¡Q���6a+e�Q��Hת��IX2v� ��$ؔ���f0��ڥIv��Ń�o��7X ����s0z7]0�����򝝃�9�ux�������k�[^����q抁ß�+���*׬"f�!�f��\�I�%�w�fr����Y-%��4���~��X�����)���Y��5��~�*
���rbqꖚ��W�M�b�d�
%6��m�Ȓ�C����J�m��B�4zU�L!�>�<��@�O@��C��>u.L�� <@�ș�G놊S��ѻ�����b����@��4��f����H�G��k��L���$���}����-*o]�w���Þ��S��!��{>&<����3kz���l���7��NE�<�x�H�MuU<>.�|;�0�WN��7��u�m~ɟ��[p�:��$T
�~9:����.O�%L�i���C�͍.�R��j��P�/�i�lE.�i�z�um��k���nU-R��;�;�b��ͳ��6<�Bh�'�L�C?�+����W^ſ%tdT��h"WeхR�ʎ����<;��"P60q[����$ngv����	N1���݋���J���
=���i?�U(_N�'��O궬A	�p�1��J�ķ�����D|K�����5S�J�������<~bz��p8<�؞%6��_ux�U#��mi*�l��Qs�����n̸�}�N��M� #�¥�'2Pg���ʙݎ��^��L�	�HZ�p��n�7E5R�$�ja05�c>,��sE+Ĳ���()c��í�{3���@�E�g�X+��y�S�Q�9�zlbi������� �9��� _�I���\#�ע���k��f�䛱!�A��΀
�i�b���wΥ�({��gմBmo;h��Fs_X���g�?>n�N����s�ľ{}�� 8bP���6��p[�h�ᔄ-�����+WMoܤ����G<�����"H�gIK'};2�ԕ�P�����~�ۙ
<�a��yO�.����i�I�p�he�#N��X�S�W@S$�FZy�;�?]�i.�QK���9�X� :2B���v�g�����~i�M�WN��m�[f���G��&���	���:j���<��]�Pn�S'�Ϥ�8>��4�O�tw��㾡�*�m(yv�f)�g�'��C�bӗ�0Ϡ,fuu����Z��� >�&[�
�"�JE������b���t[\v�M�l;.I�o�i�n�G���rt��t4��\G�	�14�i�?�&�9��1p���|o�a=~��`F�*���I����6������ǳ����L��=Aˈ����כ�"�^�H�]��QtTũ�Y���H�4��-� [�1;B��L%)99%��aT�M��:MM��C^�r�`�)8LsƔ+\�E����3?U�4�h��
��9�a8��
re���|�p�*E)����̺��-�����T��|�:w !���G�&��b(��+g�nz�Ɖo�7�Z�3^��K�����ΛQ��w^�H�^ ,i���I�)vᓏ/UYX�(ضy�uЀ�.��?��z���P��>����sRk�H�����WNZ�-��[���#�%����:��57��2~�N@��~�?Ƅ�+�
>i����RV�R^���'�Z$�Ή/w��>p�'0`�}P�p??k(����R095^�����ķC;Q���r�3��Ց5A��A�rDñ�z�O��KE%��e.�Ik�3�v ��khB�x}������(g|�0&(]�l(�u�-��@�]����|a�4������7�pͥo� ;Ӽ�Ӣ|A��a�������{w��s<|��{%4i����U���b��)Ta%H���-�ބ=��2ʙ U�d;���M��-�My#�	#��8�@�B�5Nm�v��"B:��o��Ȁ�=3���r%���)f����@^��94�f�l�ᅘN����5��mR��`+��E@E��"�cW�C@|Zi�R���JK��n���o+�"�����ke��M��Y�k�r�HR�&-_�Ih������NYm~6��6�2��Z@9Ҙ�㬑���bf����tX�ēK ��_����n��}c��3@��+�\Y+=�2��3n=������w���u���
�%w6�X�wn�c���L�1+��
,v�7̾���Z�p��5�`�u_e͙ym�ޘ:�ߤ��}QbA��$��28�~�S���7���M��uk�������č��4�N�l�-5pE��Gv���	en4�Gw�O�8�0q�۲6��|e�ǕE�̀���c��7��.�������QI�TB*S��F>�h�SBM�����GB�SN�*�|��pS��G4�D���N����S��a�0`��-8I`^�)�������ˊ��h�Q Ŗ��Sn����1���D�
��1S��W�נG�+bG��m{P�YC��Kq�P~�(�o��������Ͷ�ʳ�&���5��k�ќ�E�7Ͱ��52i_K~��V'!�0ߖs�"4�*��$�4�X�;�V���GU�Wb�J�V���)�g
�?|���ȃQ�_�L��jtHjG��7�=�s���N�O��<�3A��!Y�;4�):��q�G�C��hJ۶&�*;��HAF�*B�g+,�gh#��p�{ԀI���ŕ�t	X^��a꽸MA��[��2 ���&�$>@G�03#���`φ�97�FFH륀��:�[��\l��/��~��+~Â��z���3���XL�:~[	k�N�:�d�]=��O^h��žjY�f�<��eh.��N@ڣu�8�M̪�{[]<|d�1rw�B���u���SѶ2nUt<y��n��3��P�<n���[П�B,����M��{K?�N���U�2��YvE�|����}��qg�����e��K�������:G$|���5FAc��(E�^$�`�qܑ��WBE�ѨH�T  ��t�p��� mE�x�p��\�^&;I3��{����4�4y��u G��0��n����|Q��9Ř����E�B���ݷ.��b�X������=x� �qK�N�䨨��2&�8+��Jc�!���'��+^[k���L�H|:�%^2Ƹ��(�����p��?�i��5G ��TKg�:5��MFz�����;��������B�eݪ�M5��;v��Ղ�.S+�É�#�P��J��̘o�<�l�@Z'��]��ޤ�8YV�����}���u�v��k"403Ù�#�� ��?u��F��8�^��M�����K����|]/��B+��z�1C�{�lxPG��� a[�����Վ��LOIW�I����K����A��7�W��^Sʊ�� 9�W�l�����w���ɖR=��]�� N7ϛug�՘���	���"�>�EU�"w�7�X�,���^ϊ��)�丈o-��<�%�\�A�L�1��p�W,0����	Q齋eM�>�g�Ypn��o7 ����Xx&��^��Ǎ�Ry-s�:ڎ����&B�L3��i��o�9H�1�v#M��"��!��䌳���g�y�,*����K�$����C?��O�xl9��gXA.�.������CN4��5}�5H��k�cd�k+
i�`"M�ܔ(��3��߻���ʞ1�ؒ�Wac��8�A,���s���i[u���, nV�8�e��;�[]�}dD�ݮ߬��< ��;:,޻!>cTE!:T>~i.dk�!�?}����:2�jdd�w���ȏ6-߉H����=�a%��*θ�\�H�� ��Љs2�G\��:㐳�4
�2�4q�</��ᥬ`A�F���������?�]cv��̱
.h�bN��_���D�O��������H@2EBZb8��U$�6�	@E^`	�f�`�b�n�Y��D�vR�;0;�����C��l��!�R�m&�Eö�un_�lcW\�ڀ�*�윐̄ݺ��M���2��509���P�a�c��\�s�9��%ot�� ���Y���]0�rߑ����hIzN��u��O�"�F��Y?,u�j��C'�ѽƠ���k�y�'F�
f�z�T�~
VY�pa�7q~���f�9���z��ݼ%�_��MBvh�_v��Y2��fa �Ph4oA3랝� �T�F���1�^�΁0�l����	+�|<gUÞǜ���HC��Y�(�����b���&��`N�k�ƇG
n��|m��i�A%wݣ���1�^��w��J�ֲ���M����l+ʤ`x�<�C��5y�?�ԭ)�A�x��Lb�@Z��(�/�q�:[��-����������9S(VUX����n�J5��p��n"%Sȃ��J@�����,T�"��&� ���e��j@̸x�g���������މ����f4(�0��^��v"j���E�[�D��%���u'M&1v(<B��/�l�6�x�]-�rtW��Tw��:�� }k�c�麽��i�Zsa|U>&����MK�I�HoЫ �eK�[	QUrG�y�Gw�gOXOI��O+�%�c�X�!�� ��|M��ݜ��lg���2C��h�鿷�C�ڐ��dF�2+�̛v�7
��1��Z{Xj.�m&����ŝ7CVNLi9�H���袗{��0O�ԫ�����ʔ/���p�����z2c΍t�q�Iw��ʤmB����JT{d��}	�&���o=�#�᪍�d����H�"��e9�����k�V#���T����
+�X�oc8�����3[bW�c����9�7�Qq���5i��=1q�3��K(TԖ��Sl2�^��W-L�Bt�;���H�YJ2c�y�߳p��#[k��	�#�m$�8�j�G���׹x0#|� ����-�Mך���X�?���0`���Z�f}o�
pU��l���5al�y���xQX����}�?�(��qf*3K�ѕlNbK�g�H�%���ѵr�W�~��tM?�2sv4����T�o������K�㟪�#k�W��o��'����EOa��_=�����o7�)�Q&&x�o8��2�̪Tcn9�Mq�w�x��Yf������(��������艔9�mƗ:73�dݝrR^q$�q���|�����p>��ϸm� �A�}�]S9���Qŷ�Z�y��O�� dN_�֢���S��������E!O���/#e�x��]tv�[��`gP<=���9ߏ�SѠ����-*E�5*n��%X� M���2}�۰�G���]��[�d�䦹U*{���q�x�ʆ�T"�Wh�;?��g;N�1�Z��zd�T��h�M2{+T����}�5,<[V�M-Z|�sY۪].%��b�$s�7�J���,đ�ĩ�Q�Ռd�Q������j(C����̄��ҡ^�Eܭ�(2�l���`���xN��{���'P�ըa�Cx�Jb0����N��a�����w��s/��E(��R�	�zLq�
��{tC}�ER�{���n'B{�"��y�lVn~Q�JvĬ�#hH�I�Y�4�Ր��\�'j��b���h�-����y�� |	H&+x��w �'��cZ����g$t�����*�Ǝ̹�$) ��fmrP��=870�#� 8g�C9a�D�C-'�Y��3�� T��jγ����������b�w�����1�Zn��o����ioS�~[w����r��@��3�R)��2¸�hW��1�Ȟ�H4@ZW�V���rf�i4��������Ǘ:ߌ��/�d��@�5��zZ���<Sp��Xx�K2ch3���?�m"/hH��·�G�yrj�DΊ����=3q�BxU�$G"���B�xp�Sح�<��;���IN8L�pk*w��m�R0$I\����-y?��Ǿ��Bk����h�y�9�	%�n�[�A�j�}�H�<���)�����hk�>g���M~��W�b��9ղ�kaO>�1�<� ��WQH.��l�
�+'|��nMO�������idM3��@�MG���h�3З9oo��hr��k*B��SF:��G�����=�T�$V<��Lݗ�t�-֜����8��:����?*�ƹET~�.��s��$92���n}驪G�`x�$Sr�Y���#~`�ⲉ�$�>F���"Yg�zY����w7.���m3���і�#�\X{i���QZ�n1����@u�uaB������PC��	�i�&k��O0�K��=V��v�K�c���В��ʏ"�S3@i)3������^�z�������-�@�{|���T�?ۃfX�@��d�I��nȏ�  Y�>[��A-m3�h:�K{u�fTOo���K��a��W��axE@_����v�*݄A���]�c�G( �j�ϸ�w�bt�Y��:��Q I�5%��Ƌ��Z�aԌ|TS�w4��3*�����})�e?��=2�ޏ��[��YV�ho�>sg��.�^9�'g1&{�O+.z�y��[߁_X�Q���(��21����!Ҧ`���q��c�p��F��c�����Ϋ#��W��\i&|=�v�{ C�4�+{���%�]�-��O����jB\�:���Q��y�&�h�~���o����(I�*8e��b#!�q��=M���~��U&n������*��=�V_�2���C港 ^[��U���1b�xIl5��O��,�pt����e���&ΧS��pIt����Q ��)�䴠g�'�_���!D��E�y�ՔEµA)�r��X�q��ǽ�5*j�<��Fu�+NՔ��)T~��.ʖ���\����=�ӵ��-����wdm��UIG���o��%\.�s��*+��_�LN��&q�@����Ъ
��b	z9J5�ӕ$��V�'Z��?D���,��6(����" bR����=�< ���$�M��c�B=
�9[���p&]�&j�9>&��)��у�,�;F��Å�v��j��B��$�̬����D�c
�C�tw�(���]9�;��Mp�ao�UDd��>A1V�h�>�-��O��}�umH�?�M�.��M��9�4�<�T<繦65+[��^F�J�<_b\��F������y�%��F��^�Х�D�Ϥ��.�.L�sc���Tg5���������\{	��D@}��ʺ 8ߢt�i ��3�ѫ?��o�Y��{D6�VEI�X�i�d�\??:ͬݱv���E4+ct�kRF�7����ao�uQ�7L��"����ؽA[W�SE�&��c^�Z�!��_�Y�3�����?�S͐V���Ͻ�D5���/R��왉G��������A� qKb��a��&)�Ҥ�z�On�������b�[m"�K�)�q!�Ư�e/�5|vCW+�1_3���r'�aF�UI��9�ɪ���x �C Qf�Ji��Cz.�祈l���Џ����[:~��JL}���lJ�WY���0?��.��S�pЊ&��<[�a�}�P��%�C�ve���6����K�X�ܤ���5l��eM��A��#2��Ģ����MYz�PF�W��Pfi#rK��� *���Ƞ�&)Z�Pm�*�"Fr ����R`M��Zq2�pn���r� �!��#7���*G㷌��H�0�y�00��H�'����!�ϽP�4�#_xt��ּ�˶W����P�!	z��U?��q�)����nT����0�������X�s3lC� o�*�%N~���7d�Rg!,z�ù�\��D7�e�����zj&�dӣ�˪�G�컸Y��̔l���V.�P��|�����Z�0���|�f�H9� ��=
_�$�#=���#o9H�V�{E��)5,!.Ņ�c���9iƹ�\p�l�ޫ�H��@qpKE������'Z���h��I������ ��v��]�g �Z�`"�p�q�pځ� ��&��&nA�8 �ԟ�j�Mc�0nI�`�ozϻ4u��}(�.M.�ӭ��K�F���M�I��᥁�j��h��Ee٘"��Vz��6?}V�F��@�YI��O����qQ�	�eN���Rb�<0iz��n��������u��+�)��*�6���{ȼ�o����M!�-��3�����\Z�Xa�v��n~����=�+M�2���a�����XZE>��e�EVHw�v>G���������������pP��������7�� ��sP�����PT�de�MrFE{��m�6����� ��Z�J����zE�Õro�P��K�����{c�ͽ��DQ�՝�n��UG��V�\A�3b���Ԯ��/:����Z#HUN��"�f�b'O͎���KÅ��`a._T=N�Ϧ?��J���	s�ݞ5�b=س��F�j�J��E4�v�A[;U4��+Y��#�N@�%�V���T�fF<���@��S�EH�l��@�	��kߘ�a��#���vb��
�j���!o� SW��������}�Q�C$��CV����h�E�p���-H��2�>�T�p&��1K���㷚�xv�XQb= �+6<OOZP�֦���(#x�R�¨������^��
X��%���!]�*�/j�7�'Q%)5iE'�l�͘#�n��)[�#���M{ %.���>�$�Tb4��4)mw�exPQ�������&)��(K�ԉf��{0s�3�?	!Hz��Q2Ua��;��݁tuU�&՜������7��\�c�~��y�cS/W�?�u�X����WG�e�T`����iW���+��G�Q��Erq�۴�$�^P�������z�Sc,l}\Su�����B�j[S�m��L�Ȝ�ֿ��w��i��H��<�g�T��A�@���Ҳ���.Y��@%OSL���[� ��8�[���6������ ��Vƫ3���3���bY�PiS������)/�Ki�n�<�(��fJ��s��R��4��]�K�K9�]�ȵ)����IВ����Y�y#�,�{��S�(W&U�4*j~�ޫH��D�zM�翎���&Z�IN�)������αkx���>唕z�UC��Z�z�BaO���CϤ�$�-�
b�o�Pk��p��5�a�{A:��yl�	~'{�������,�W���ƴ�0�p�����K�[���N�ѕvy�deW0���HR����a{������VcD������dA��+�a���+t���:�E���>%=�k����^�z"u�m��ɢ�D��BHv��А�7Uc���sD3�n!n�b�|jq���� ���|3�_����&�lNεq{���w&j�B�Cٽ�B7�I����_�5竷EȪWp�JG6T�v�m/CA�U�sB*!�ͬ@�#I UT����N�U�(rd����@>�"�X�Qfc��	mpQ-�����|F��5��$��:���;<�f>Euk���Ĝ��X`"�Z|���N1s`��-=�%[-�V�.H�M���\�\[$�U(0jP >zK[8i1��C�L�F��&�O�J6�i=����@b���� �۵mB0�B4��|@$�є#Fn�aW��o��A�g\���g���Ng������C�����qe�j�w�v��?є�HHZ��xTo@2��4�wk�S5��S�> @�&�����;bﾲ��o��3�uT���Ѯ�bT;H�$if���5�Q��a����1g]�� ��P-˨�Y4kgڭ;3̔o[�4�e˰��$P&8�jI�qC�����;��d0��&��bR�n�q�Ĉ8�h������\���C`3bk0mC�/��վxZ��>��3����d&[��ו�_����䭗 Lx� ���58
&��_�Kى�{�W_?�t=f �%00�^�oVA��T×!$ؾ�[�ȺN���Rjy�y�]k�}j���P�ba��u��į��~S�1N�Z����_J#
+Jl�of�l�Z�Dx���r�@[9����5�6��w��P�n�P�������������~�*K0?D��Yu�"�dN�����bd�i���PD�!��~=�ts~�O�3q�e��Ui������/1}��aTR��,i��t,��Jp]�F�U�1e�Ii�h��yxY�.�������-� �Ĳl�B�0���>ʟ�j:�dV��x� &mZ2�K�@3���ܢ�v~�k9�m�rB|�1�a�DV@(��i�H8��D�0��tۉ���h���9h��&an��ta�t
��p�b����v6@�&�l�5?�����I��5��j��t;��Zf��봴9���w�i�Ӊ��݉�(��͋/�Ջ��f*�|����)�ˋ>}��bfck�E��U,F��(u��$�6�`�����A�)�\ٱ�2�E�U�L�-����  P��;*5���h���F�x����xo���C$�����Ze�?��js�:c�%����pS2�������f�e�}R=*$�I�A�_&Py#g�T(J0��E�hu"V����,��iu^V\}��7?���!HAf�ZL�[h:�����F
�~���* {�z��_���j����xj��B�`4s�-.kNΟ�3Z!_99��������hV���R��Na��}D���Z(�|c�z�V,�|d�)nX�V�"���`&�l�]����WVA7����'a:q�B&u���K�0I��2�cr��í/�Y�+%@!)i3�MP���ab?�t��t�����!q��W"�k�=y���k��6�񁪾�1�|�x�a�h�-C#���}��uL��D0�D8C0P�u��?߁���"��Tv�Iml��A��^��	�~J��:�:���	�Ν2�ԾΎ�h�5ozD����j�V��?�8̉:�B��Պ�!�
�a	�^���~t�3�C��p &��6VnT�c�(mO	����y+q�cʮ�Ggf�o5Ñ�J�Fd�܆\]a�A��Xj�8J#K$��f�^
L��u�� �.�W�/[�ݥ7���g����g���������@(�(	����ߊ�C�5�4����.n�a�/�#F��<�ˑ�D�X2���JA]�(��p�\�f���Hܳ�%���qD���8��)Neo3_�5�6�E><��E�c��$D�D*/\*_�A���^��,K,;��L��ji�JJ�d�`���7���uӒ9���4�Su�b  0�2u�&�����k��U8��sQ��-T3�Яv�^Y�����!C�}�*ɩ
����b-�iQ��9�7X!]�$ObY�Kk�$�#/��JONz����FQ�\�Z�o��~e4�{d��3�(�"y��ø�
���L��+L~�9�$+W�\����V�w%�:t�C �nY,a��z��mx">���A��4 j�W�l�`�B��*�̿���� hs�U�'S�T�:�J�jG���s%G�NCZJ�
��A�����[�����\�۲C nZ�&�|X�}�.P�rE��b�o�u�O��cwJy��x���Pb�(�%&�h@�'����9ct	F���rmg�%.����[E��C��񇊷��b��9��U歂��<��
}Ҏ.�꒵�S!�����H�J:r�hh|-"G���B���H�:Q�l�#������
&5��Z���3 �C\�y�Z̖QQ�����U~��.��]�l��3z[�;g^!��ϫ���,���_aV��$��i���ص��kV�	PiR&�������}�'�j�|�����&ˉC"i{��ߪ0�̨;!���Ũ��0X=/����'��|1���f�:<�v�X�_�^,:@7~n�� =�"�����A ��͓�.��>E�C%�����L繁�W$C)~1�
W�bU���\=i��K���jQL[0� �	��5��=��H�B(���P��y��tJ�fE����,E�,^OJW�%mՙ�x�L��R߄��A+#l����_���!����g�,u#�w74���k	���W��=k��H�\�7��:M��x]
8�gr#�#�����A��jw2�~�qd]�k��{(1�\ui
�xtp�GQ��(�/C5X�k��7�eK�� {}��M翀]�礡n�z�/��=z?��^���MK
7�pWPwH��g�@��є��$~�\�e�=�4x��d:��e���� l���'�#J�nh�S��U��{�ِ~��+����)~t�(�!���l�����}�V�CA��N�K |�7��o��4�)j:T�q��k�s��P��L��f��"FM�-��B 7�㴱�'���d��9��o��g�����qYG����dSPv��$Y����+a����4�xك��e ���6Z�_&��g���On\�u�Ik!�&~p4E��CN�s仯ȉ:Zo �fT̥�Vw�UOp���Ht�� �\�� �{������#�%�L���υ��f5�&y[Hd^y��?X
2=m�m��bl�wy3
n��V �0���RE6PG����j�gO��.,�`V���*�߷I���q!Wѐ��j�B��%SQ2k�mM̏/�!�W	g��D$�`�����+����;�tw�jVhGhv�'f�/��l�s��8sՂ(7�L��-�\���\r20���g��95��%^e��ɧ��h{���^|$�7��J����6���[�߅�x�a1SѴ*�B���]��Rɦ��QI����'=�-#D�����ѧYx�m��㩺v�}�<�WI���.�����C}^���|���ݠ��&�1@5��7�"�̕�=I�'І��ϗ�r3�)d���(�L�<k�E��ʲ��d��3��gdNY+�N��A����Q��`U7��M��Z@��^Ձ���t7V��d<WU����dֳ���1W�"X\S`�ű�&�>փ7���q�A}�Q!٧���4��}n��h���h�Y+ 0~F�_��+�mA9���{���ftb#%� �xE��;� �'��x~�|�@\���0�*E�j����#�b�5�i�u��x��ZE��@Y�!�)Co ���;��^(%�aQ��*�V��)c9��^ �b~�~A.��̦5M>T���_�U��*�n�vc0�6֦�i��'
��n`�%�N�׶��*L^�$R��uH �uȴ���E^?�&��Y���_"�Ȳ?#��ςGl_l�8�D$��-ZrfL��6�h�{�g.
�O��A���T��| k�᭳��¾֔C?\����/�i�
��d�0��k[�[�������/v�	SeH[V/U&�T�7Bn&��;G�'����&`����%��ùf$틱��4��+L�\8�W�qzav�1�����z��]�����6X���ȡ�O���3?w&w%vɖ�kV�B�k���B�k7;�R�^߯���)���e��O,�6A����E�
���J/��U`Yf��d9�8�u{�I+
p����M#�.���d���z���Hy���ۅ���{0S!q�2��/}��������vn�H������ANr.c^�,�t�v!����龇U2�y�7���N:�4����膛R7z�*g���"b ���@��+�آr��6���E(����'���ɣg*Q$�ڻ�`]|t��Ap��6����t�~	������x��Hs��[N��.�������
�3"@t�M�!k���ϐ �nq���j��Jw h�sMj���m�;A�Zrv��l=�������\�th�E�Ғ�tΣ�l�B���]���D�?:����sD7suĲ��,�#�Ha��r��$l�%���Zrx���x��ǯEy��Ko�p�b���L�P�����=�!2�![�P]J�g��#5��/p�_�Z+��j��o���k�֓��^��z�v�[��jK%
IG���3��|]>���$%O��Ԙ����.0.�h�:c�4�G�44��_�2���C`B��u�A��'��ٲ��d�8��S'�̰���tr�Q��`Hʞ�MJ8�o���;�?�Nc����d&���NdwcS���GUq�wʈ>�&_�c?���G�c�W��+��AJ�ո6Ĝ��&us�2?*�n�7�N@=�.׷C��]S��xhY�8) !`�1zU�E��}>2d�N��V�tm�|�yVU"GS����Y]-�8/�$��Ԧ�U�\s>r�L�7FΫ��A̜�mu�𪆭M��y}���as�q�HȇК��c�K�#���o���,����J����r0o�:5xG��{<-�����ʡ�`��;��&X˃�h��0_�BY��Q Qi|	��Ggn'mkL��T撧D�x�ܾ�r���������]���!�#�[ڄF\��q_<^�^�hU9�`��<�����o�J�q�~�:"�Um{g����������whojF�d�8��;}�Y�MЯ:�V�eC���={S�-��s`����V��
�AW|�xk��n�M�D竃��c��� <�W��X��1�����]T�Y��?��z^����å��RŸ�_֢Q�O�f6�;�Cf�Me����)7C�f�=g���y�� G:��%<;�^�z�E糧I�� ��Q؁��������d�|��?](��P��z�pJ�<��&|n 2�؟����zұg
�u����bv�G�5�m��_,[(��}�E	؝搜DØ��_f*UÌ�R��ɲ�U�QNA�NV��2㉐���K�3�H�?����J73�;[d����=��֔k�r��JD8�s�j��`mľ�˿�-�Տ8m����;a�äV*v8S��/fj��(�4�x�8m��,s�e���T���3Hs�����-�AH0��D\"!Z{ Z+�̙�#�����/e��G���)��j����R�m��~��I�>݅�NABH�tR���=� �	O�A��q"fF���5�����N�7�>1�q�o�J���~ŌwO/m�}�1�M���n=
Q��덚 u�m��t��3.�bݤ��#l��*�S����iو60���>�~N�'':x}���*��!�P$�<y���Pś�G�'nF�i�T_e�~;2_m�� ��rr�6�΄>��"v4��ţ�j��\-�=e3|�^�U��u�N�8H�9�}�_:JFy*
@�5"d�H�E��M�V�1������$~�^d�Qz�^*3y>}�^ijX@��� �'�{�,���)$��}�O.�f���\�:�,))�� %�&��2��A+��N�M��vm-.Qm����Z��3��.V�ep�횝���q��k�l�y�j&D�3�� @�$C�׺7������k׫��v��U�g�6�x��ך:s˞殆#������CPt�ʔ�C��'��k^��sT���l\X�R˯h�+���>F�K���H#�nO��7���;�ja^3��/�?���Euo�+Tg��߂�M�'�ɽ~��6h=���x��W�ԌxJ�3�f�997����&�`V���Z�����?�ٵ�>�Py����ZP����N�{��j,�A��Vy��cB��~#�B��@T�4	:�6��,��a�dx�8o7w��m��ž�2��T�u�UϦN��ʗ��"�R�c��NR��(��"CB�~�,P��x�'�vl�o ����!�����C�q��qk�%���y�)�-?����]4�O« L�>Ě@�Rj02^�@piԫ"y����E�3f���^c%�9p����&�Z	�����i��Y4�o-�T���B�~��W�_ӧMT�V�T�n'@+��lg��2E���d��2	��n�gK��^&XZNx~��6�s2�ш��mIĹj�U	69�1��X�N��ϳiT�&��w�`��j{�ƨ	��|6 o} %]?�����%�ɮ(= �������OOs�֜��G�lm#��3[�C#9��iSJ)��?��1����r�Ű��Ç��{\���q�)����7h%�)6��u!^��4������0̝��4�D�2�m�d�րsg���R���L�"�6�o��_c�Ŭ2A����l�T��r�%�W�)������a�x��ǋM�5,%�I�i{s�,���2Lit�����P� �_�0���a8#��w���1TI�`\���Ъu��a�n0z��}��OI�BQ�vE�r���e;T��B��ïl���k��z���㬖����-���gn��LK��Z
���j=oo�c��2
5�w����g������$tw�砒�&$��4L~v�}q��5X���F���'"��u���"T�)��\G'��8��%��槉I�}�JJ�W��F��;x�Ģq���J�@�X	
����͝�; �昗��ڍ�i�	�D7?�LN/0$h�C����Cy�5�_�aH���WoZ�;(��=��pE�r�,aFNrĞq%Gp���3)ǖ��U�����GE���Rl���l������h�a
-D%��nB*�P���&�����l��X4)��m��B�9=�W��Wg���%y>�!�*^w;�o�Ъ���!1[e�M<Rr��mѐ�kA�w,�J��'4�j��[r�ӯ�cz_v�l}+�8:��
�a��z�,ܼ����ٛ�:��M�H��\�Ӟש���Jl-�ʸ=�E��N(�Mc��C�U����)&H��?��������HkV'd�5|K�NGе��^V',�oO',�1_/k
��P�g�)�<���sbPO/i|1�&:�J�%Z��|�#&�����2�09�9�I��ѧ#�л���8^z�M/��������J���5ky$
N�Du�W��0����1,5�θ�k�w��;%���Y�-v�&审�Ee+��I9s�n�j	�G�����F�W���wrh+�|������ϲ�x�QVv��u��0\�=vD��-��̉#�%��CQ������C*3����+�@#����G3���}�f�XU8ww9��H��j��R&��RRU��݌Q*UQ+��i�#��Y�bo)����O�֬��� KU���+N7�jZG�[#{��h�Xt���!z�I;�v��>���
9l���W�3�FM��X�k8|�ru�םU9�ȩ�l[�:󃘞@�����0Ao)!d�3�,֚*���k��ӯ�1��ad��8V�p$���d�B�v�ob��U�ʍ0�4vKܚ+(x�Gjݧg��.��_mF ��3Gx����>ҚB�2SY������p"�/�"��;�,����7��|�e+̲�KQ�rO�Vw5���&x8�(׿g즔=,��-i��Ҝ8�\-�m�v5߻��f���|a_�&�޹K�I3�IO��\H9R�v\��󪇜�1Q
�Bp�<���3� P�����.jK#�z�XT�v�W��R���L7,�"���s�u��M�R;҇�����Ê7
��i�q�|#ܫG���&��	��z&C2���y�{e�`Y�ωjd�2��2HY��J�����jL!q+�MN��h�;3�� ��`���ْXzS��T&#��}0h�����\�9I�4�T���4ŉ]����4�����2�U~"�SCZ��N�s��J�l�.�u��l
�1�\����`e� F1>�c��Ƚ&�44sI�D��X�/�1o7��^C�O`�q�cJ�o ��0�͏c�d�s�u��ej�w�'D&�8�ܲ�K�N���(Έm��<��;=ڣ��N.�=L1��x�(\��t �T����ZJM�x�d��&d����*�Ni@#U���w��x��L�~G����'�G3���<jz�1c��稬��L��fW,&l d�Nؤ�=|�"��a����-�-n�'�䧁,�wӼ�̇(�ɒ8B_tJG0��gԋ����ܦzGo��A5���nx7	S��/�2 ��֟/xm��%)/���a��ބ�yٸ�+����0a���t��$��1�����8�OL���d����'���p��v�ʪ��2Qzn]�y8Cէ׌�a>w�ū�*y�F�X������"����z�e�>�WA2%�����1�˘䉔������Z۲v�;[�yH�J��kQn;˯*>��)*����Ȼ:̘,�G�=���h52g��n�XBI�� ̽�*���Vb�-�:}&�1����m�U	�Ȕ5g��p�]���;�a�$��]�~.\�a{-���y�H�Uhl\7n�G�*�`���;H��Ӧ�2(��Vå~������w�}N��)��
�O]1��2?���j�[�y�S���4qT�F��%��Ϭ�g}���H��l
P��D��ސ,��?��4D�G�`7��	.B�ʬ����p��5��:���_�	C��t1�	t"*?V������&�I��)a��Ľ����^\3����˗��CC$3k��G�U*�0��G㯈��m3-\	4>P�־֡�0Ób���Ļ�ýu��L��"�쪕e3���&�(����j�/�
�r
>ş�iT��A�9"w��"Po9S��T��b[̲EY�ݿ[��H�G�P;ݻ[l"�=J5j��bB@6���Gٲ�$.����G@��A�cQ�@�7HG�#fR��V���Q�u��#?8���kxe>q�����A:M���;�E�����d�C�kU��y���H�ԍg΍�`��]�������9�ɲ9,�0f-�X�J��P�����ԑa�#x$��slc��bnm��]��괫 dR7?��%��JP�ވ�K�{�`������~ퟬ�����0��Z4���S)��?�����կS ����/$4�;��	��,���dK�n�?�\&��P���˒��$1�>����61�`)��7�7檈�qM�h��ڨd�{�������L�}�p+t�e{��Dtl9����p���K��?��t���;5��o�-MEo��by�\	)��?Fإ}��&�m���/Oc�Cs��2����Oc���N1�q?�تEoB��h��j/�����8�6�`�p�MyF-:�Tc&ӫ7N�����0)�_ߐydzwp
�FrEu���o�dL}��/ţ�{�������wоC�>��d
���ω�޴t�޺�}��@����b���٨�4&b2�����,4�Ir�p�8����V��,��D�ou6�o4�o���X�)tؿ]��@�����;N��`B�%۟��КpU=���>��_}a���/`Ńd����uy��^!��}�\�F�0�r�3��5������}v<�V�Γ���$��'ȶ�p�$���M�jV?"o62�ʁv5,>Z�(�$c�v>7���8`��1ݣ�������;����� &�}i*NӴ�H�$$�ќ��e��F�kzǴĉ�ߊ� .�$��N[6a��/�5k�p�Q���Z1	|��\��1�f\G���D��,� >��X�맥q ��ϵ��<<o���but�<ơ&��0m�E����T�"be�<���T�"p�;ӫ�@�6��e����^��o���)ãM�����J��޷�S�P��U����=^�����c7ż���˦:�i'b;:I\��HVՄ����?���s�@��hQ"��?�0@�%���d+�2Lܺ�56��;�aLs��aV�S�"ɰ�D�1T�?����=�{I�t��z�F����$5F��Z]�$���h�*ӕ��P+��G�PE�{\ݭ&k��x�
-�+A0<���V�+�g$�������GP���ܱ���n���珌������}��W��bn�X�ߓ��E��P_�N)Ϲ��r(2�g�C1[C>�����e�G��k�H�"'�����s�h���� �$���)LUv��1#E�5���3�6~��x�*�>y����v�SA��Ib�K�����gȲ�j�)�N�Wm��Q?F�T�.���y9�j���Ն%��hA�;�e�\r{����F��n���[���wMJ�ry�R�E%�O�_���큁����0�1g���Rf�W�a�u��r��>�&�� Zo_�_D��%`�ޣFd:/�w��K\�a����f��;�L���P�n�5�������.F*�v��V�X]���v���W[h�m��K�!7�g.��
�2�u��]�j[�+P��i~w��|�!���m6����T�3l����	:]'_p�侒b �HJ\T}J����M�����
�cb&�tS5�/�F~��Y�΃A�q��L��������x��Rp��xՕ��1�#�~�ME��e�2�k�ٯ�����G�O�?�~�~2i���#��W�@�^��%؇Q��PZz���R E�vE���{���ʫ'�iC��Sr��<��VZ⁪,̀�_�$��]zăw"Z���H�����~do,	-�p��fv8`wM3˯����!S���N9�ϰ�Cs^�H֟�\H�?�\���k�ƣ�3b��eU�vﶒޯ\ӖY�{)���R�����.f��ɴU�G�P��G8��R����.d�żf��.��v�/���fh&D_�}�9�:����붹�ހߍ�3��=��-�UJ��]Q��5�	ZH|��=�A� ?�Gh���B�8�`V��D�u*�(�J�ׅ
s�~����H�uvU��\��L	�`I�/�����!�A ��~�-�ru\���ǌ<�~�J�_c ���7v�-�W�Oܟj_C�:3ʾwt��(<'(��DE��%�ݫ�|w���fT�}c ��'�����x�GԗR��{��p�����]�������ȷa|h��4��j8E�@�)�緗�����x�m��xѯ\��LL��̾|ޏ>�U�[�*��ƨ�\��z��Ci�������8j�A	Oq ��|`���y����V���ۄjI�6.��d��X�9�ֻߌ����ל���]������6��e���Ii^;�!��.��C��+Ao���N��T�0Xi���E�A�ў@�^��%AB�o�I?}F�֦���S��@�Ҏ$�W��;u~�#����"r�р�o�����Np���\��em8\m����(3�=��RO��70�MU����K$�;��� �����oڍ�61(~02h
B�݌݊�UU��n�8A�g�V�mUPo�=����{m��M�V�e`Q\��us���83E̲ݯ���K��S�Uf��R�~����Ճ�����=�T�P�+҂��&���~���^UuǬG��T@�@���^�?i
�Qʗ�������ֈ��I�&o!�p�*[�0�Ѳ� �xdСح���Zٙ�Ո8����6��%�� �5!��K��Niz8��Y�{��/*�3]RT7�?:��i��|�:�j�))Ѓ��A��{s>Ю� ������.)ByF&�p�kW<Ў�hy�V菶� ^��,�
}���i�!+�g=$����Sg�:Aؼ��l���\'����/֛��a��&>��=�]��M��H���r5D��c/MVF�Ν��b�]~K�L��͜��g���<�
Y^놖�gT�d�!{&��BM�W�8/P�iՐ�a�������J�%wҎ���Տ�g��l{��A%�t�M���0�te%�~�%����.F������,�T�~���D��� ��kЮN�Kg�St�'�oӷwM5|�aHg�i-�}xp��+��M0jDo�ȱ���v�E����z��Z�3֥��n��T�=e���N[�ck���)b6�f���d����,F&�L��4~�o�(��V���1*���+���&l)N�C��='G�+�"F�g�q�*.�&M�f���+a��<��#����C�,6��b��	4t�х���+x��òڀ���5�f=}R��t|���P�{�xEʈ�л�X�}��p��:����|pLQ���i���P���t�1���Q>��'t"�,o�p�%�p�[�5����{����H_o5W!�����e'
-ȝL�x�V�<�������y&�*\"����X�ѣsF�R;՜<m�0����A�
����FY1�D�����%>s��,/y@��\���e;Tg�El7� �"��õ��A��#A��̉g�t�Gt.����5G�f�܆�ncOf�@nk&�����\�^6 ?2�� �lh��deO�m��G��6}��1�3 Y�:K�@���,��v��I;�0E.	W��$F�P�\����(0���O�����g��GRC���i��0s�]l���4J�	��T7���
u�V��t<�j^wl��5+2���]�SU��AՇ�y�K�;���L��V�w��u���P�s�����uf�u���I��Jf�Ղ�9�c}(N��x��m�4���O�{O�{�jg3��'E4\8�������栻0T���;�R�w>�ካ��0"@���_c&��T�ש�O#˧ݦ4�q�f�4�|5�.�1���舡E���*-��6d�H++��ϵ;W�^�E���[�����?H�c�$�\v2)I�SOB�p�E+��ݑ|���ʼ�2�>N��Ct�ލr��P�C����9�"�(��f-Z*0�c���U>:=X���s��)L�p��ɧ��"���T� �WJ��N[�}t���c�ާQnq[yqܽI�{<���k�k~�?ѐ˗��h��ٍ݅��U6NR���Q�Ybv_��#�@�*S�)�1��q�ʋ5�I��v�rӫ��x�����=TD��$�X$1��[���L�&�y����5"P3�z7�$�K��#)�p昽*��g2n���m�DM��*���"Qfߏ�ĥX8\'N��b�;P��oi�	��f�}�!z�'L�oug��-ۻ� ��5�[�a���k�^ڌ
��������W���+c���̾J��0��6]�f�Vl�'���^_�2>�WE��r77m��b��}㘔=u��&�:~�`���7ȼ��9�qo��r�dN�=8Y��	6OcV󛉗7=�����Yx��E%l��6O�n��w�~L5���r����D��a��������A:m��������r��gv�F�aF����3J�s<%nI�P.�C�b�TH{�����e�c'�jӝ�m�sʁ�bhM�ۊ�9�y[i2��]��L�jG���\�Ֆ��y�X�A�!K�,��D�>���ۿ����_їm�Ի�7!wf���^Ȉ'��S��N�t;0���{���Q�C=�ǟ��x��
�30Q�r|Kd�7����CO �Q�>%������@�_��6#q��K��4�{Ah_ݹ���^ױ��P�~27�/�[��vv�gR��Wˣ���H��A����l^a��$I`�"���#���88��G��m�
�\��6��|�պA{C�R��~:�)8���ǔ�a�7�"/�;�'(@T5�7лf�Z4\~���=B��;Ks��`.g��T='�����b����W$W�F��g*��Ѻ�c�.� I�(�ر�W���Oؽ�Z9�"����$��s�����u$�֞��E'�����=�F})3?)�`mvz�!�l�
_A��%=M���qF���sQ8?;`�ӈ��d����[ԡb^���q�i����0�HV������ɬ'����^�H�}���8��T�� L�����	> 
m���ߣ1�׫�f7� r��J
�v�ӗX�W�s��\�rs�t>UJg��T���ۥ2�U-�9���ί��%5�W�Y1w�R;�}�[X��Lt�"�OG�5���>2"H�ӊ��]i��@��<2���"�Ű���@0�OJV��&
-������i`�����A��u	0l\��Ґ2A���}���a���DWKy� E��;��M����$�d���C��iH��SlHCL3�4��m�1ua!�B�=�z�5�Ȟ�F�[�1'���;�3�.	tb4|F(�J#����`�@���z�"5�ﴸ�Z�8f��y�ҿ�e$bw|����Fa�)�:��wan}l���mUOl�Q�]f>�[
Z��F�~Q�2��)2?��VR	���&�zOu��A���~c"�B� ��#������nK2��*9@�������9U�S�&d9��k�9��w$���n�<b0Q�e ���!�5h�<�9tK|=�b���:ۂ���6�i�t�r��S����L`�F�]Փ� ��p���]�Lu��@�M_���^���P�.��B�Z�4�ix<|��:�@�E�6a�������?A1�t��.n79���N��WQ@��Xkʑ�+7�T��kV����W�Sj�j��~�I%��D���+OQQ��ȯ���e��j,��,fF���ãOIαE���]���ewm?#�$22�uT�cmIi������ȗ�L�軦)׾r��ɚ"�
�h4Ғws��u�z�|ɕ0����)�GP�ۺ��?B�=�a�,�u���"є������[��ra�Rn ������LCD���)v�;���Q��z�w�K��Ԟ
������i. z	g]!ƈl\��y
�3v�g���iE;C�T��,s����~���D�/�u���Ӊ4l�
u`'9]S�����&x|ڀ|JZe�#
��X�C2���`��S���W��d.\�NpɁKɈ^�U{�Cc�4���rw?4�ݶ���X�h~�l��9����G,	p��-��P����b�<.���c����q�-�p��bq�#��}��N�φ�C�w�`� |��M~-�Er=I�#Y=yh�pțxT�I�0�D���G�t)}0����k?��t�~U�9yN�M��8���f�Y�w�e �pK�o�L*xUb�Џ�o��O���?�Gh���-�M��J{��9�}��/>R3���!BB� �G�J�Ӈ���0��O��52�F\�1XDy�P�麯��v��/�hG P|����5��< ̏a>t�K���
w��܎J�&C���<ũ��:ݘ�*�8,�wd�(�g]g���8q�ص��Η�N[�Q���$�M����w�a ; �d}O�Mg��`��5~���D<�����qŗ�g{��1�������N�?�c�j�_��������I�A2�<�5�[/ҙ�ٚ.6�}�k���`�/ �6b�,<q�ϴ�
����0� _7�� �؏f��[���YV,j�t1��t�{�HW��`�W+�ef�ƫ;�f&^�=A
���MX��~��̃�q��s�Ɔ�S�O�m�7��J@?���ն�u���[s�]�WW����T��	w/��1�Rh�p����� f��+C��X��K��i�n&	]�L��6�J⛣��j�5K+k����]
F�*����6��"k�nz�I�c�W�_�B�G�.�y?޸}���m�TP�JJ뾞�/A�/QW�8��zW����W#l�ZTPP��ƥ(iI��b�% Z=.{|;i�#�ѓ_I���]�L���R<�g��_�{�v��t)=�vB��F��,�I6=��I���NhY�W�5w��(��z���X~��$D�	#@�;%����f���u��rg=���.]6�j�v���ĕ`e�׿_��0����@{>�o �/�E�H�"m���Z��Z��F31?���(�O7Z������C���U�'_:L����O���0ȧ@��L	�_��0q zS/o�$U{��E�cr��d���+{���}�.�ӎ��#���V2w^�F�w�n5����2ֽe�~jB�m>�Vt����!d�C,�T��@��G������ ��z��Y]�Sc[��n��GS�����C��$b���C%�N��A��6��Q�����1�1�[�?{�Έ�g��Ï��AzQLk�����Z2}����U⚞j� 'Q�M�&,(IH��߽��["8��� �
��i��>��ӟ]Y�������CP�t{�"��Ӕy�2?�N_�KZ6e\�g<�"�ǃ pb�]�lj�J���8M'��8���\�����#���/~*��ߊ3���ax���KvDϯ:�������/�/���W���\��`��A�ջ)I� �����C����JҚ�+���Ѿ���<��i��aH����͞��1�Y��X�jݣ��`ƤZ&�I�/ME�*fJ�N	�G�g$@�5R��x�z�r���~&��gx�l	��h,`���""u���#�
���\�*���tr/ �(��>M��g����o�v=���u��i5-WW�7k���e���u�F�I��gIe�Q����W������+��LC�;��c�/�`E�-��C��x�2'Y;g�3E]Q��x��^u�FR�3�cRqv=�-K%�z}L�v9��X&�i�a�ʺ��&���x,e{����*PLӳ7�S��Yh�t�H�T��L���y\2%W������������΍��Rrr\I�zYH�Q��9f'�c`J��:=%���^G�&\<8=��I�s���W��'�Vji����c�s �_��o�\��M��B�$G��+�Ȝ�\��(�E��]���q���4�z�t^�V9��������>�,�%7!��w�.QW�{���?�uV2�=����m+ᬱ�G�!���>�RhO!5׳ZL�S��Pb�R�R�6p�ǎ��`<�"z@V~�щ������e��b_;��?��8%�{l����Q10+��a�2#F~�C��g�28���if?��ޢ�#�d?L�Xe3M/%6�h�^�֩�f����-�|!2�<�����8�}=����T��K�Pb�4��z�"�X���B����+��;2���a�=�z��,5֘D�9=_O�p�6�P`O(cd�Z,��{�ƬR��p�ϒQ��<��1��et�C�q�]�,k:Bu���xT|6L�&�����%s1�BD��+�%��6?�@l�c�*�E`���l�ש,~׉�!���}�j�c�v��mVs��#��1A������Kw���US �J.��u�/�ӡB;=��C��9�M5+xoB�l�\����z����s6�\Lv��͚�L���'|�Y��7�0s�
�9c���nV79{w�HC���� Q,P]e��+ڂ���(�aVcd�5�5����[�cA�% 7����".��!���%�L[��bXWG�7�vʂ]�!�{/��,����z�֘Y�e�b�ly�Lz�
�fim|\�n��d���?�����,��rg���|���#�^�_�9�_����D����^ )8cBC��߫�8x��<���eFPs
T��y,�KF�OM�(D$����r��C���85�K��3Ŧ��MUN�al@����=��j�������aLZ�^�7�NP�⼘�]m�P=�'w��a���Z����is�����}���&=�)�0��q$^�K]s��R@D�8sc�P��h�hYi����^cm%~�}:���K�t� q/j~�2�Љ���9�T����sg��"P �{�����m�^j'���Z(o����n��W�w�7+��j�.��n?5�C�aƗ'�2;b��P����\��֨t�QN	�u��u5��~��C�w.=I�|Mڨ�
�=��s�����Q�O�(���2|]�[@�\���Ƿ�\s4F>F��-�0��dm���[����
�<j��&.NKy���&���$�K��RT �0q���	f�$4��/:������a�e'�h]��Rw�ǻ�� � �Đ���MVז��������Y��zS�RdW��)@��6[��b �{)�p�D���5zK��2�#06�8�~�[�:/�NoM�F�0ȩ<����D�;_Vjϫ	 �����&�A������(�n��b�%:v��!��x{��˅�RW6�,!�C=�u�I��q�ه�D��Q�K��D�r�a���h�A���xMc�ڞ=Ⱦ��H^/[�yTϱ�V�O�d���'�@�m٣r����\�喁�/���$c�� ��[b��>�a%{��I�9{"�Bu6���.ũ֒��J�kK�(؃� ң��p�KZ���M#�D�b�������a�?Hu���e_�"<�z��̻��$�2}<'2W�:Q�7�ԕ�i.�:+�:	���%�^��K�_C���)b	=�<����ևw�h&�2����l����i-�7L�3����ոR;*]�y�������j?�0+٠�&D�nK�������F��G�B��S?kc���]�" ZseXa����4j�=��� Y����0���K1�~���ec��>���+b�G�ɉpqߨ����4��J�ȋ���&�N�G�aV�U��}~z@��K8��QIt@S��G6��XE��ρ%|D��~�b��;��|�m�����h�t�`�5"�H���p�!X��S�94���_�=�u��\	�c�����&��$y��j�!�bB*�b&���2����$%�ow�dr*���(�[�}��K��=O�aE����ak����L�M"���vU�N�1�ґ[`��::q�%�9f�#���g硺���:=Z��4�����А�/p�ТG3)��F�.lhA��\c=��S2��X��',����\p����bs�F�A�#���Y?Ї�tT�0�Qશ�tv-s�L��0���i��:�I[T��,�]A��2��C����g��-	L,�	��,��֠]J�j���Y|Y���T޲�ӱp�~CF�%?�Xm�4kL�0���E�]q�aOR��%G�{�J5A2��˦�AG=RھaAi�]���X�B� /\Ž��3�xb��2=�^��DN�,�	~fC���]�) ��ڢi��>�$U��6�v݃U�
1l���[Q�x�<CY�b��
9G�*J��c"t�lQ���Y�#�:���ӻ2DG�KL��C��e�yiK�#��<m�t����P��`�bʶ�$.�sF��Ĝ �'���d7�n�ݎ��pL���U]����*���5�jl���2�Gl[.aH^,vꮛ3�?��6&�ؿ&IM�ٚ_I��x�ꞍД�lm{v`v�p���$F��c��?w8|(ul\@���#�yκR�T��<p!���O�7Gȏ�����%�c}zK����N�T���D.=&�f+�>R�h�g�h,_r�~;����,�`�~T����M� ��lb���w��\��=��V����mY�Ixtr韕$��g��i�I9��L8�E�lS��k�	'�)���ڌ��AW�S'a��:��d���g���wgH� �{ƺo�W�P�nX�ß�%s�j�[�d2�����(�u��5֣G!��ܦ�֨��p�>�N|M�;��l���/���x�D6mlU�����?���c�{�2E�+���	�8�6â���������P�Ǻ:����a��_��%�ų�z2Vre��U?�f���6q=oM��0�j�4�̲8�^sӥo$z\�!���el���.�q	#����; �Խ�Q�3����� V.�dH�^JB�-d���6��R�P֨'E�4hM��șܦ�Z�|�a�I'>�,�t_�
^ɘP�u�h|�V�;&�	f\\�L+�ָ�Ʈ�#1{�Sr��T�&5n�Jz����,_2������N~ސ7�b�j�H�l��06AD��Ÿd^Y<��L�@���A�u�
ϒ��� ��*�ٓ� J�}� ?�,h,�ʧR���b�g�c�v�e��;w�*���f	gV�-��(���Z;�L3����}l��D$_g�K8i~ݳ]T�{�s��GQd�$�����O��ӞF~Jc-�-mu�D?�5�3�B�B�ֱ.��ιH<�����g��z���}�'��;�gB�����9�bK�����7�{�K�WePy��?{j�^�ѷA��D�����=�\�S}�E�SW-P2��������b�י8�'yM����m���R�v���]�R�����x�vRϘi�&��oW���69�p���������b�&]SX��76��M
�2^�ϝ�Xm,�D�~.�!�E����i �/R�n�J.�-��(��	3Ǯ�j/B~�	���1�X)�oRmJ�	���[m�Jf�d#�7���;���I
L�ֿT���V��;����۞����DR7%G�D�t��	�	A�����Ft�{B=4� [��+]���k}�8ĵ�͕'s+n��|�PC0���"n�>^�70N���h�%P 5��խP��	�B _��cd��^}���%0rb��U��6!)RcPNVM�0��v�ȡuUM���'<��
C�w��@��s���ٳhaVF%n��&;o�jЕ�W��w�G.0x������� �P������3�.fܠ^��g�F���K9�� ��؞����Y.�*%�A�5ه$R��R��
��[��6 |d�UT,q���t;�%�k��D�{��1�s���'O0ct�I?�7���}@�ÂE��M�^5̆2|���EZ!�&v��i"�"w��@�V�x�?ջc�7ʬ�U����a) ���N��6<�5`��DG����I��ᄓ� ��J�6=}<J�?݁��9���1�)S����ra#V�����j��1�0�?�]G�����<TC�0�Q���"P��uS7F�R�wP�
�8���g��T~)N[ti�/�JZ��#QFq_.�n�:�] ����� ��U�H��/�ܐ�wU.Sr���}�m���R�>��l����K����޾{��n��:��b�qd�K��߲AM�,�{��H�0>
z�`�p+%��+^\� ���3�[z��$=E��)Y�z�y�X}�%���^��KRes�غ�����f/�)_g��K^��	#g�SϜ>]��L�@�ᐮ��>"��nb �F���b��p-��J�L��*���l�]�Vk�]��%	�g�(��:�xg���v���1���X�\�e�{^JIy�|�Zo��gBM9�ude'a���镅���0�C��a�t��$X(9��+7&��"�veD���4��;��[�0&��{�_^M��؊�Ʉ�L�=�K��TJT�P��ܛ�ug!����(أ�(�]窺=[�~��$��I�`#�~�A��������ϱ��`��Uc��k�*_�&�������{u�WԦ���z���s+`���)��"���	]�r}P4����<���7�fn���P� `���
|��c�Du?>`cw�#"B��w�S�����7�zϑR\Uf�~S#�� �$�ܐӊA�!T{��<�1�H��ƃ��a���0@�ޥ��r���Q�Vy�QkJ'j�1���#ֻ񇱾�@�� �yRn���B�B��j�Q>��+���y��K��8+�}�^�T�ŧ�,�ۢ�~g���\8���\-��4�?^��=X����{�����`m!��4��bEmx���8��:�z*Q��gy���+Շ.���m�wltM
D&�f^��	"��l`8_*�T��'�]S2��� �_� ���lɘQyڒj/�A��u6@8�&�H|DO��{�9�n����+���5�E��|����^����@�
mb��Ӷ$�`�q���r��N�h�8"Vïy������=߷����8�i���L0B66�S�=�$ ���z4h�o���d�7��Ԫz�ʨ�� -cM��,��9��[[}u���P�:2$�h�a���%�j�e]����ᲹeX�_ʪ�!8���G����N\�P"7�#!�DJM�0�g?��o���*
�6o&YI:m�����ج �gI�#�y`��0����$ú��+d7���)�� FHƼ�#��B
R���FR�~�'"��%-@��4-�c���Ѓ�����.pY��Λ�\4UC/V�O�TE�8ϗX�#�ؖ���B��6s�\�?N�����w�,�t��wڬ����|�z�eҠ����Z�e��u�7�򡓑����qj۽�����������o��@��]%0��
�41�W
�jwA?�AIp��\��[��Z2�ZWԻ&/�ˍ��$�;dM��rUe�r���v5�^��5r�˪fA��t�q����ř�ȃt�R�������.zJWʻrM21�X�L�9��{�c���#g�)ɗ�f�����C�'?k�=�C�:��g�8��1{��S
�7`�֧C�Cr� jgӓA=��F<L�4������J8�����Q�3#�4�{����SQ�y_��i���r�N��B�#��ݲv�����9�q������V?!닍�m��{v?0�J|�`#�;w6P�U�q|QC�ٺ��k��cQ�B ��!]�h�
�%�@�ł�Ĺ��¯����~u"JPTz<z*��#U�����q�E�= ����h6�G�́���Kh'�/>�a\��=�L�C��@�������6�CڐS-y�M{�,��x�DF�_A�l���[yj۱K���h�v��"FO)�s��L.}+���֋����BL�o� q>\& ����_5<�0�ENϬ�+�
h5M�(��@��g���:V,�x>g��D�N���	@K�+�_�l.�S�h� ��~��epl�/��6} ��X�]8�3�Zi��՗S����!���i#�cf�G�s#\
tn�s�J*'Ζ�n�<{�x��м�t��oD�7R���(U��#���?��*s�ۼ�e�"�8n���ж��Dm[�)��1@+-%�1{3**$R��`x�,��D.!㡼k�QEu��3�	2`���1M�WJT^�iFū�a~#Gne~�F�Ĺ�C�܄��0]Yw�3C�a�몃��rȓ��qŞ��j��!ǗHp�5� �9�9����7��Չ|�ܶ+`B���ܧ{�� ��(H5�V#e�e�!�3�=�oϢ�\��E&L��g����沧&��s�h�|��O���5O�kp'�1w�X�~��cl������]"���M/S^׽c������wn֭�_)#��ɵa���7j5Q��l�4k��۾˾�,Bt~������a����}�N�-{�������1#��풘��*Ì��kcj�KS���d��G=O<؃t���U܀����J0�<�PR0�[J��}��9}-�`�^S���]b,�KԢ0�����ь�8�đ� ,չ��Z���@C�H��f�ۗD�����D	^Foق�
�p�����[�����zIM��Y���؊9�o��W�qH<7M7����B�.� Qb��,j�*O�(z����u�|%/y��7�Ht�u�EQ�\����'��}�%X��Ǯ�o�Ϣ��������� ��k�:n:�퀠�dqB-W�~���~�\mZ�s��Nr� ���7��p�+�5µ��#z� �?�DӧƗ�fi8������]�y|��u������u�rasw�t�t�q�� ���e���6w(�0B�E��'��C�F����rh�2��.�[�,ڹŸ��v����_m������h,g��swdt���1���m�x6H;2��g����fs�<5�r�u�^�v���|5�e�e��ᮮ�����9��-\����3D`��\�����o��j��5�7WS�%~b�&�#��z�)ϓ��]�l!4��0yA���y߇���V��x%.L��$��K�Y���.@1-S�׃��T�]����=����#�˳��t�V�>0\��t�a�k�4R�9��|����&�����F�%�8&j ��9n6�@	�������㋼���~*��4%�ԥS�*� �.� ��De8���!s�U��f��Ol:�.����[c&��]��3����]!�/5{����G��M��'��Z%s62;^���u�XZ5
K.��m�_:?l5�Z�ít[y�?q��KW���á_�K
����W?�M'F���fj��.�{�8W/g�9+Gx��r��\��ɘ�m=����3�X\����O�b
�l_[�>�g8a��t�����,ă��ıB�������6��89���g�ɗ�--�T��*���/�X��$�~Q�\'u�ЁC���W^2�*�	+B�j����L��hg�:Ś�;����p�(R�� �0�])J������)�	U�E��r��1@�ݵZ��M��sd�[��DI�`����s�:�@hS M�w�Ŀ���24_iߐg<���g6�)�KEL���ڲ��)i��/�
nGh��-~��5
y7�t6��>/��/dg��|z!oC;K�t&������d$$"��G��བ5���g`��0�E�LJ�lw�^��'Ȏ ��S+��ߥ;��u�v���Ҕ�[qc5�f4�~��� -t{ᯨ;S��Z�Ss�UCy�����@B��n:f�F��D��w˹�>����.���78������|�=��o����u�wjS
˾���I*��Վ��yV�n��Y�Q�#�\�6
�;��򃾡�h���F��|'��S��(�1IR�D�I#��}г�[�U.��#��6�8�^�c�)ۯak�]�S�4�-ނ��MvȎbN$���S~�}~��:�H��z��u��勻fd��T�'�&���U�R�0AH����GR�h�`b��|f�mh�r�l�~���"�Z)s��-e�o\<Ӿ�p���?w���*�M,{3q�1�ꀂn�s�N�����d�x�A8>�|$gt�N��V��6~�5:m����r2nUSF���m^��v�n��`w����X�TtVWB�^-K��7��u5�gHMپ{��F��m��q��F�A������a�M����iX�]v�<%��f�y̎�2
P8Vh�����|-�.M�ɕ��(�f�EG}]N�w�X!�E(d�-
��#�;Msɖ�cW��;�/�c��1iN��AV�a�r��N#�PJ��v&'2��Ӟ|"��Οȯ��8( ��Xг(��Z�dκ�è��`@$GEF�/KA{����]i{dnKB[G��Db�w<�(
�$�[@ؒ��VΛ�(M�FSؗ�;��8�J�I��"d����aS˨�qʠ�\���r��3�����,6���7<A����Z�^���ت��+�a�T\ς+�@H��x�eR��J)��JBA��Q�}F^�&o�5�����Rf�ǃ��L�������M�&�>���B��2~�I�)�Z���@��K�o��{#1���}�y��kq���C���tŸ�B����7�=xou�8
a�H̝Hq�d����IB��l����"I�\={k��p@�v}�X�� Q���Pr�уd���b��ɝ���=��^�ʁ��������$ ������.":�?��oDQ5���J�m���vM��࿟d6l��(����M�q\��d�3D_�N��)�����WN�����Ж4�|����f;�x���Ķ:�tB0U��/����i2Έ�%ǅ�ȷ���!qgUt:Ƥ֊�=�[�����;�⺳�d�A��5�8�i�xT����KZ����� >f�!,J[jf�Q�Ta
�F.lӎT�X���vք�n�MOmZ�¸iB{����`u��_^qE���eX�vE{C���;0"�]p\͙jB�V��PQ��6��5VRpv�l��(�S���J{qUlw��M���.�|���z�SkO��G���B�1���	�l~^�і�&`�3G�u�bGħ��%h��/��"'l9 ��i%�ضū�P�k���ʣ��\�(T�t�ŝ���Iz�B�Ձ{iX@[F|������>��34Tn��q|ZT,�P]7�S{��w��/ހ���.��DS�8Q���˟��g��F�si����=
{w���>A�9����"8�f�nW�_U��� �!�b��-��ѧ��3I�GQ��b^�α�e���8J0�̠U�>�|`��Q
��/���(*�J�-p^����KxR]$�IP)�_(��^��
d�����;"�$ş�)�f �!�-���٤����c�=(=Ϝ��kU���y~�b�|�w�2p=�QP�5��c�A����(K(��w������[z�������1��r�6��7�����q3�9.w�%9�E8��Rش�"�k:�@�p�W��T'���g���I��F�����MĄ;╷3(�$2LH#r@G�������ǵ���q�,��-�]�3:sW�!Y�Q�;a�����o�ӮH}v
���B�?�rI����!o��W	3�@c2�YG�R�?&���$yL���PJ�Fc!�lXzPQ~ڵ�)e�X���j˞�b
ΌcVs��ix���mq�c[7Exj�R���KcVLvvU��XJ�c2�{v�5����f�D�$u��׵���?՞�m�F,�'�}9]��q_���[O.;�5�:-ZG����u�F���H�cEC��3�s��� ����@^n�g����N'$�%Kښ�ن[ZF������/�qHAW�3���<
��)��=1Gs<��e�p��
���`ks�7�>�/��R�;�+-�������+�O��������Þ-�����H��æ{��i)Q�H(Ͳ�lL��
��2����M�ͷ�_�	m���5[ḣmOd[T��>'R���̘Ml�e�V�3�������*��
S���,�׃z���<x�MXC���2;�9��A��'iDS&T�̦W�����[�b[������_��
&vԆ��3gp��Tfd��%Y���ꨥև6&�{�h��^`(jjC<#����W��S�3�[u����i�=E�d��#�%�B�oS�L�O���p�1@�
���l��|n=+Ã=�v�2�a�Q�� �r�+�^x.y������H9��7����ɧ>���\��.��_7E�u,�u�/r���C֣��p��`��+��ާ�����.�T���u�h�d&�^�T6\l�H&�6:M�z�!3+Q����n^�v���Ҽ���((����6b~@Y��W��o[i���	߃�pͳR���W�����ŋě2)�(�x+4rC�����V���Z;)��AىK"y-=h��Dd�p@�1���8g�iY:fm+��F�A��}��g�1W�:c:ǝK��1�4Ƽ5�YV����/@W���>��_�7����
��4`3�Oց�n�2�9�	��8�׮F����d��f?���V�U�����	�@�
��͵�����V�C*�C�ʐԼ��Zaf#�Q׶�Ҫ{է������������⯶�"5�Wo�糚RQ�4��h��r!#R���2�OS(C�b�ǻ����رm���v��T�Ձ�V��Rl?���6�	�+��6��F���ǒ+�:��Ch��fo+�V�6��~�CdY��v�ſ��1Ԓ���M/8w�#�c��<�b�$+k���gR�(����dA��r��dr���� ��$`�.����l�=,�޶���Y�}BD��3b�0��2��t6$�24S��&A�b[�>�t7�&Q�s��w�8��u�HfH]��Ѓ�J}��Búy
d�~�k�\�p��㻢�o�Ej#�K,��>m��S�2zuF�3{�}N!�JB]�UHP�f��0�$�͏f��M�J�����g�<� �~E�CB�N�9I�}��,��e&��[+��������{װS��P�jp{��q���ל�޻�O���^d�Hv�� J^�u)�~�K_�!��k�At���e<�S�ml\ގF�r��ޜ¬�%��� ;cbr��g��i��%v�y�����n�*�嗑������Ń��a��M�Ͻr�5P�_~1��zR�>�<��۔�$�����lxd��+��=���#i�����M�q�4�2$�"DDS��b��Zh��~Of�LY�����F���o��K4�������Z^���p�h�|4����7+�Ӌ�G�.��6(�9Xƀ�{�pa�;s�o�:7g%�B��ᔧ��;w�����g(�Xh�����[�r��]�u�
��~����z˔X����{�;���H���ji�����U�,�!,<<B<}�;qzK��H��kܨx�p�:�
\�g��9'D`a�ֱi���~:�@�&���)��!���hϾ�_%�:5� �����1�[x>0s�U�SX����B�_(���yV�l�/a}9�k����,�ŷUB .��X����;-�C=;p=�np=X�Q�ט��M��C1ɡ�Й#t�i.L�g�@� ��7zP�?^-p���#��>���n��c^e�;�;M~y2_=A*�	$\.���U�+��k�!ع�S{�9���6Byy8�2��I����O!��U��ĖA~��5 �
y�����%���AV��:W鹪��(��*�E ��!>��G#���Mu���[PgЅ�#�aM�X�!6����.��)�n]WFm�A�0z��34�#솼%��:����}$���n�w����(�tE���֗�u,������p�D'�M�XYl��0��,�I����<��]L�D*5魗�JaE@3 ��h�ql=�e��	b7c>��rOw�P���GG0a�)S.�|���n��ퟘ�x������j��c�����[�a�,cO:�Q��9z�>���ȥ���`x9�;~KU�z`K�Zs'�"
^�=�Ae'1粱�� ow���޾T�VQ����rZ�!2�r������%�̺�<]ܞ�����q��7� '�1��E:�����6�w�7��\j���ޙ�$��)11��T����!���x+�4�eA�(ҏqy҄�#;Է����k>;[��A��V����7ܢJ�K!ҚD�����#%��5�^��^?8
�V!E1��-��lQ3}Ԍ���0�q��G��)7C����	jɪQ�ˣ8�1�������K%��,�2��c��;��-���۲3Q)Ū��p$tF��TF9)FV����b�}�o��ؗ%FǸ���8�#q�g��ޔ>l���&�ꀤ������D���.Ä��k�(n�z����@��j�D�ż=!�LH�Y*�'�i�N<A�O%��6�C~�EGk*b.�7vap5���!L��"»9��G��{�0:E���!G^����-����H���<MM�,�Y%��茔a��_��G'OP��eD��A���!����hPƨd�E��:�ŝ�ܩa9����������a9��d�˖D�wrurX�anϏR�6���|��O�XrA�0����� �<ٺ��RC�U�����t��w�j8�_./+ݍ�N|؆�Ȯ�^����S����6\V����0�rr��o{ʚ�Λ޼�C�J3��'��n��Z��Nn�>�`NS5���7��n5�7�a��-�47X�s���b#0��:�~�"ñֆK�������I���P�C��A���~ >�����IfX�Z(�G��dQ��#����v��q�-a`c;¿]�&�C>?E;"��$5-�
v��V�ub%"Y:\�� �17<����늘��ݥ�;)��5l^�C�3���(�YX��'���|��$���WϿi��Ef�e�,r9T�4���
Ʃ�t0B�F뼧��0p�l�]����u/����07�I�W���a��߉����(���!;����u�oU�d3gG[2{:%�i�2�(�
.i�����`2k��o��vEWH�ܻ�e>����P�Isz��N��:���(��w�B�lZ��=���F�p�Z�m�� ���S6��C�f���J�z�Kͺ4Xl�)�Ί[\G9�d�%z�Ӈt.�� �!ڍ�H��W
����בap
o��A�i��w��jOH�_�u��c�D�;�Q�����w���L���K���)�6�^�>�`�:��2fZ�Q1s7�����QX�
T$�D��9݃~-7H�/����/'Ze�Q�Y^�G�j�����m�aWOV��\���Cz�x h8����b�^F;����̜��/�R��M�5��`�&�DQZ�#v�
A�5�����b��n(�����[��p� Z�(]�I��X��-BS�{y~e��4$ \��v�*ي�*�la.?�������!O=�UInG����U�ZQR��:�hT�Vi*��@�]uL3d�A��B����S��HҘ�T��n�H@ƫ�դ	P�%�P�MZK���v��I�ڢ7O�EV�[�;
��+��{7'�i�`��ZP�Nh�6nbC�;��:zEXC�sͷ�ŚƻW����s�>�JD��qM.��c]Ҏ�E���-���E�;���+#��A���V����^
��"6��`k2	�Z�%h���!X�-�L�y�f��G��R}7�s2#Pf}���x2���m�AF��
���.�os�U�Cr�ݨ±:�o�sH�4����ʭh;v�|?�:�
I$��Km_���P��h�����
x�p����k���@���xo�򗹘�7�|�����ס�,.șj��'hJ�f>>�\27ov;�9�;3�6�r����j,4��e]�0����_�O��2G�yo���|]�bJ����jN�f�א������%��I�"Ҁkr'��o�b��q�!6�VPKk'��;?�s"���;�U�WQ]�l��ϡ�e�h�^(��{�֮��U̿���,!�j���z�3���R��q]��61�zCDN.��{��I!�J�t���A�A�k��=/�EA�$���_K�6r���֟B&��S�-�!�UG���yQD8~���;OS��'ֳlCr�D;�S}�@eVʄ����~:��L�÷���u�T�g����Yor�����"�XV�`0/}�h��-�7�������g4��hBx�G<e���s��Pu���=�fڀ�+���O)L�1��4vD�i@���U5Z�IR���I���w�DF����J2��Ό9Pm{��1�Uy+�e��K�^��TQo��]�yr%9��|�A��L	�YSI�'z���g��X�@�K�H�#��>̖�0CU9EZђ�	$��)�Ò���]�H-I,֋XCđ���@8/�Ϣ^���g����;��b�2���in	�B���4�>����ɹ(�[�h���>���z��o�ݬ������Ϲ8{��ޝ���X��,zƭ���"�����|s�4�X�0]��جO`�4�8X��W���E�S�]��"���\��O�з4pm���z�^���6��_�]tj�`�x<�ONF�\��
J<�Y$�];���9�ak�S/8�S�PB75Ot\��>�c���;<�$�d��.� ����Vk�O�%������T;�6c�]F���k��[�)H����;��SlSd��e�7g%g(�A�>��'g�Ęb!(����%x,+j9�J���p��x�R��&��d��F����Nj�K{�k�k�n�|)j,m�66���0���$
��n_���A��X�O͂3��q'2Q4�%zG�eN �p�&ӊad�e%j�*.$Vbu�lR����(A��.�q����i�V��<9�+i�4�>s���;�ו��B:^ލ�95��}ODCn�pl�O��]:����?w�W.��	���ԋ�VC��70��LY�>���V귯�"fL�~�x�	"����h�T1 ]i.>[�E�K�m?�=����DM����� �Bώ�^�|�Zɣ�@������[ڴ��R�QTc���ܧj`�ZQ�?��sa �k|H���Vw����.\��?���G�,�K���K�Z���C��*�$��{���D���4ά�����Pr�*������LyG�}��`׃k�i���k���͘e�^�:p�N��z;�"/g�*�h����_����; ��Co�c������O���G��xoG��e�Ү��^��з:��aٸKp�� �í�� ���
vCg�̈́�^ػ]�Y	�_1������C�F���d�\�R}��7�m)��1��Ҳ3�_��~9lk�e!��EW���~�P�]?���.gQ�$�aW�Q��y��w�'��G�?~J�S�%c<��Va��q>j�;����>/r>��2U��(Mwѹ�g�%6��dj\b��3,��M�S�T�eP�ۏ�|9UV����n__�^�%vR�2'�;H�K��Iɞ{�Q��j蝦�9��2�)��b?p�%~%<������L�2mj��vߑ��}�7�D����V�B�˛�*`z���oKPY_�5Wpjn�܀�n�P �|p_��K�?
�, !m�B1��� �E2��4�'	R��W>����Ң�J0�k��H��j�L+4�G��Ʈ��p$b먋W��%�KCk�@�޲W��'਴5��VZJƞ>Evr����F1InL�!8��t��-���(0w2���~�{g�%���D⚉K�����6����O��������GKGJ�\�
�|�D�j��y�Ϯ��v��hf��x�i�]J��i�-�G8�����6����]���XdC�)hmI����햒��8kR�	J�q���$�ɘTC�mh�掽ܫ�ǉ�'���+U��Ƈ3��Ѱ	y6IGd�ʰ����,���.;��2����2������$~c����R�b%.6��� �a7m4�(�O4/�%5K�x�Le��!+̩rq�>��)�s��&87�1��#�@�+������+G�R_%��(b��l�9���Hfz��D���y��Y�g�Bh�������؆8tX�uS��|A�x��)�\�v���^s��lC.D��#ɫ�C�Z!.���nUW�%������D'ź6��h�A�^���
B�GB�� ��c��.Y	O㥩�������|G|�C���fTb{�~���4�<�r���2}`T�>�(��F�yx��R�_�4�E�*;��xdӓSb�f?z��v��ˎF�Au��ʒd<W	TF�j3�:l�놶:�v�ަ<��C�pu��ѳ����@�=��Ԭ�0T>��B��y�2d�M��XC��~��^�����́��\��vD1�^x0Pd�6�1x�I�A��*p���e��k���Y���I>]��Ru���5iOb�	ϟ�D�E8�}m�2���M*�(��������ݜ�ܚh�������6�p��9�Xޕ��@�����] ��s�����O�- �pP1�-a3˧��f�v+gذ�Kkܟ��Kr���n0��Ya��3I�Z�k��s�k7{��o�Z`:U��l�IӔ�NJ��~�XWƀ�ѕN���M'��ѣǎW�����f��,����r����pv��N��_`E���c� .�gھ�Ӑ�7�Q48��~%���y>E�a��+��E�!��9��p[�q�g�&i�����v�2m�nt����h6A���[J ]_QU�T>m���9Ҏ��e/I
��$"d!̝�k���|rpLK-ʤ���E���oE?������� ��"���E�
�f��9z+�ʁ��~��[�j�k��z��/o�ܼ��z1�\꿾�8�o��\�b�����`�Z�m�D��$�0�W�\�����Le�4�圊֯��]�lq��/�>��i�~�S#6i>Zi�������y����+�LI�;\����E�9O8���cUp��΁p�#p�Z���M:6n����F[׎;��Rd��i�������4% {�aw�M�_��wp��t�#��eE����՞Cm1
���ީ@�Q���
���M ���l�[�>��t��o04��ei��;��S^��
����k�.<ff޺��F�g���ΐ�[2�0dF��{Ȃ{q/v����0(���ȯp�16ӫh�T�Nx�{-��X/D�	���n��@��g�Î"����ӌ"i��Ab	��S�Nd�E�<��0X��H����,s���y׿+>+�ա��=Y(VE��nlۓ�Z��>�T"v^��.���E{z�:Pr���əm�A�DD����h�^��\1�$l��=J���!�7A9����|?f���=F�i4��B�s�5^�B@�o[��C� �[��G�*�NK���
�g���Q%Ч�qA\��6b�o�������ju9�C���t����oW�����p��F}p�keE���	����7��G@�" S����r�y���w,�����S|%������b�ax���H�Sْd��_�-��e����W�1���6�%�_�����`*�Ul#�-n�^���߻�4唒�<�g��u�U]Q�{f>ͱ��`�bp�N���H��#U-���k��A�&d��)�{�2�a���fv"��XB(���h`.���/^2hc$zff�c']�v��w��t��O��MJ(;k��n�Lu8C�6MI� �!�+��{<�
�m�s=��`���π.�M(/B$��7C�Av0Y���a����_�D7���s,H����_�M�&TF��7��~�|<��
�M��:�����^���Q��_&�J&N���r���_��5���7bCy0�Y-���sG��(��K:Ǎ=���A{|n(�ΓjH�>���k��~1O���\��=E����b�G��"í�q���=�(ǘ�E����:f���I
��"�_�mU1_�����)o�F�*�c"����e������0v,�$��_t���Cx�|e�}C_ԓ����\_(I��I�\D���Hy�TR�6���VyC�Y4�\q���� �.����g{p�!�q�982©�/�,���w����XŬ�xX��Ŀ��e�����-+xhv�q������0�]+��/�O=bk��������SI�'\8Z�f�(��%�R��n�E�<�_J��� Y�;�e?%�[�?,V	LRu�p5����'��C>M׵��Ûn�Ƹ�굤b��ϸ�-��kE�!<��'Y��γ��i���|y6��ảys|�"M�Xvٮ}�	ET���5�H�	�(ۣϖ������~����^�t�M-���Ѹ���j�Y��pݩ����ώn1������>8?�<���y�IU���.{�\mz�����ʺʩҷ��q�4P6�D���"P�m���%Ґ������u�d�nPs��>� ��j^��nr����v�T�6�]�YάDi���&�G���wO|dJ
�
.��s��+զ���Br�ܓ1� ���t��k��D_�������l>�.?�l�8���rʑ@�?��]Nj�\�\�y�ް�7F��l��(��s��ِ�����%�l��u�L*♖��̰,d�r� �sv[�O �G�S5�٩JoAw5�d)'Ĝ�O��9�^Ƣ�MGV�='5�pO��88�;[t�d�ތY}����ɸ~�-�f@&2\��̾���%s���2�@ׅ��l�=5xkP=��:.��8��0���
�8
�&vM�8��9v"{0����d@��0vi��>�|�9��=�X0�(�m�p���g SG0���<�?��
4'e�Lϵ�2^V~���a����|��N��<�&�lN�v��H����U�!D^��B�5Z�Z��>��4���pNG�9T/zJ'b���ˈ��4����0�=5nԹmPmϺ%a�VY�;4;<�5����d��_�[�Et.�<5�N�a�|��Uu:���^hzܞz�7}�6�Y;��cm]Ƞ��C�����ʚ�Is�e5�I��)Z@	t���K���e��ۣ�<:����8fOyk�ϧ��\������?�!no6�'O������ܣC~��	��>) �#H_&�~\Z��62J�
a��<�3ꥡz��鮰4H��D�S�A�Y{�f�6x�I�)g����-=RVt���;:�\������}�5۞�7-6<
���ϣ�(�2�v(?3Gq/<���5�1V��t��J��p5vw��B3��@>��	��c���)�
� x�3FzV]�sh{�Z,���)�	Uх[��x���W�	�-�C*�J��>ńm�D���S�J9w�_��}y�/�ˣ(Y�{����x�a�m%�a#n�_��ݍ
_D�ْ�)+�c�À�F�fک�ߥ��H��i�8�Dp���m`�N�9A��>���{?7ͽjZ���I�K�.��(���ʷZ��*��vl{�
^��0J?ͩ�գ��5C6��=���Pu�.�vɡ#j;��&*�󀋂v2l�`��y��b�}�bV�����0��F�߾y�	����+r]p!`���ؒ"=�C���ri;������1�3NN��{V��U�ZH��laW�p6�1Z"K���i�= �˓zGH�_��DJY�KJ��V��O6�\�+��������U�$�[�1�왯YN=�oc�ն�p��j��n��(<��	EWY�Z�m�G����m{���� �Jd���Z҆]*�`�E:�I\�7��#h�bAbQ�a�9F�'�عE������ޣ�0��"��h$�����9��J�1���%�i���1\�P�y����8���F�
Y�*"�/2�b���2�ޜ�ޓs���/��H)���З��>��XXJ�`��ߦ�ڡGi���-dȤ,M\R؝5P;�M�\�V���
T��鍔7���4"��mz��fyR�y�s��k�%D�S��݋MK-Mz<��R���9*$F���O��t=!�׵�WJ
È{7^�I<��ݣ��Ӊ|�RF���N�E���՜��9�9�?�S���xB@�p�]����S�Q!�� X�D�I���j�p]g\a�����ﰻ���@�d�ɞ-+���-:��i?gx�C��Ds��T|��%\��]�����x��b����|o�q�gq83��rh��_�|z'� �9TC�NĸO�����l�7�Z�!y���p-I�D�O��K�is�<elN��ɑ���ѵ(b�ϕk����C�q���� �u�@�帎��le�mU���.�Wr��� y��뒵�ف�Lkl�i��O�i�����訥��ɾg�K�	�+�=, �O�j3��
PJA/"�+�K�C���et:�c���AX��ϣ�D��!���3�Vx�n�������b����tȁS����b��(�lEF�x[�ȇ�(��f�X�D���،���~��濡���u��6��� �m�F��
�m�D�-7:m���K�-�B?C4�^�Gc�0�e���J�Q��>�b����wy0s���A�U��[]/��}3Ԗ*�.AW�̝�ギ��ݺ���ԓ
���������E���kٮ1[`#�,�as!�Ӈ]l��^�h�W�o(ouw_�_��ڏԹ��gN��u���9*�T�)�5Rl��S?�@k����us B)�%�KɣAR��LÏP����6����ᫀ��@}s3nB5�t�P�oA�)S!ە���Mc�,c�A�ڿ�H���'u�L
U�)*��0� �n����[2�@����a*�uJMN�ԦN��M�8/�;I�?��������ڬ�¹��2��Hd���#�M������ ������� ��X�vhT��3?~Cjf�*Hu�HY�8�L������B����Id[�����(�'A�m���^��l{��qAq��&Tj�ƿ2*�qo^�Ś!"u-����A|�Ǯu�`Xp�wq8�{h�U�c{^>�k�| �&���R��
19!0N�IA+U��P���s�����iq�vDsKPͼȮ�ϰ���\���w�|K1N����=ۣ�w{ku]�ױ���d\���6��5�<��5PAE�\7Zs�B0�׮0��� ���Q���40��eGXn�B���=�GPz�����V߆QCH-��A�V��(��	p%�x��ņ�)��gPtO�#�a���"(���żȾ�����(�,`R}������ ~�3�Rd��"�9�x��`����!�'	��1�����?f��U���*�4��Hj�� �b����P���ͰF�/O{&@���l],�e6%CsF7���l��7�2"��`/w�T0b��\4��P���b���XOe��m>'*��M���54wi��b�/b�)��ir�#.<*�: �G���ov��H��i�������RR� )�<�j?dz��_����(�J��uN�5-�q��k}LSw�Y�p�+�=�~�wR�u��*���ӛXȖ+�ع
g:�Xx�7�K y�ud{��jv)ǈ�i�b�����|��x�7,����Y��H1����ZxwGT�B'��;4 �]Ta�L���d7B#s���l���eP<�83*���0�s-H�k��c�
ve��V�r�����`��[şr�Ʀ�#��~�2�����"L�(�U�ѓ�Ißj/�q�lr��GP��1!��$��"��B*�CWn�S�cS��S�(�e?��IY���qz3G��"���ݍ�75�����y��@^dy-�;�.��]�v�f�w�wz��j3�D[qG������f�r�`��ֻ{8.XV�B�M��n*A��t�
�-�9B%>0��ձԿ�|���u�>Y��Q�
�^��6=��9�j#t<bװ��F�Cd��L����Q*��L#H�5��w����^巇���B�\P�SX[�0▂F�%A������@��2(Νr�~э��|X�B	؝cR�kkS�1C���M�^��@_�����D�&T�]� X7	il�l�	{��
8��x�_EG� 0|��Ř���F�n`.G幤uo�aY��kF������vy��	m~��	E�D���X�6`���� *��@L�����P(>��fp�����bI��):�c���Ϯn�B��*�(�Jw�}'P�N��?Lp�wܧ.6T�EP\Ub�4-��&"F@&��p�Jt��ϒl����`lѤ�@j������Tv
��On�b�C��*[S-lͦ�;��Up)�x }�LŊ>�� .��ʋv����Lƅ;�ez>�w���zu;�r����^����������� ���':���A_�B��2�:"�.����w�E�n3���B�B�X�7�$�W�{TI��dwJp&މ˟��4�~�,4�����PJ- � �@A�G'ݍ�����q~+�Ŭ;,bې�>C%������}Y�1'�r:�;��JM�m[�E4L!7��J]�m@�6v;��b�Иڋn���s͕j�'�G��4<��c��5@z��L��LL=ck�[��]�0كH޺�!��t�]�o�M0q>E�l�[�vKR� %������a�N�Zd$]����yN��7
���WZKZ2w�a�H���0�U�����cgf����64�qBk,�F{BrY�x)�wo��Fڿj!v�b�ݨ8���im�3[��vޠ����n�R�W�{]/9��!��Qs�t&f����T4h+�~���<���S�%��{_�j�g_������X���2]z*cr����oQ^����=���ɘ�Zߨ�|R��Wڔ�L`�;��N�<�Sv�-}�G�3�OM@�\����e�9�&O�%��r����s[>�flc��@�-�}��E,ż}��9�ЩIh��|�S�\��}�&!��8h�1g�6*��`>"[F�96��)skˆgL#��
G�<c��:s���3���*�9jǭ}3p��R���>�+�i��a�rE�P'�c$Vx�Zñ?���ʐ�׶��H��v` K/Z�8v���.�y�+5}�_W �F��P��w�l�,A���!#�9O�aHN3��ӪG$�����J,�[	���-i%dO&4Uz���$��L��Ȟ-vg{�v㦧�א#�Iˮ���b�i�̧���~({���<e�W[�bv���v�O�4�����׭�hp/>}"�u����|���+n�4|���߳ M4n!� ��!@I��\��3�e��FR�4o�=�3)�	<���r�0�IF��VU#-{�}���t����;l�]ٌ�7=$�}ƔPð��Wt{b�<�"pYN�.^��Z㻭�vR@6"v�7��M��r��L�Gv\|i+�͐�o��Z���!X��>��1&p����\E�e7bOXD�̳:FFD�a��$����&,W0��V  �O���dm�N��[�����G��	"���e��u��Z��C��(�D�e�(����MFP7�XWbi����s�:��*�-���rZ�ĂEz^��~��Yh�� ���J�Y��(QAw�⡭�?��t�2�_k��O�?��HP�C��3z�7�\e�mWn�~|s�s|�W$��Dx
�4]��ǫ����"�7�@
����j8�x�d�e�=`~73
$�	Ы�8N�Ԟ"�U	���+b�O��Ki��F�\���"�2[��3�ټo�fN;��gM�]U�����a�u
��Z'�3�a�ـ��#	;F��cHq��.���)|]�����Z�ۙW�T��^RE��=����� O��l��OA/�1�0#{5
�fJ��`iZc�Sz?�oq�,��E�a�y/��ݪ�W�E8=��Cn�3>;��і<Q=�!�v�_��EʑP�'���1�r�	���5�A�W��"�E�ө�"��'J�H�w�q,�O}QFq:�':	�}��z�X��������[F�w��gh~[~�2 [&�8_5�5�]eǋ����YG��Ɇ	~+w�Y_3�|�M��Tɹ0��Ĥ�-��@�y���$�oن��v�&^��|4�F3Ga��u�
6��p;��{=D��C�@ެ� Ȃ�t-��[<١�n���5���J�g��N����#��&�nhΗ�#:l��] skXQU�!.:�����=���/$�kG��ǡD��?���z{g���%*�
�}�/�qїw.A�3 �n�jcO�Ԧ[���>ZO-�1�\�������3X�y��1�}Lj鐰R�T��!*Y˃c��H��\��Ut=�S�y��Ɔ���[�*�Y��9�rF��S���W��%a�4	�V�}�Kȗa�kVH �7��)��G����{��52�dL�
�I)���tV9��2�����Tw��?N@�17�3�
%+� ��!�.	���{��y��hN�ϡ6�1��@�v�j��yz� YTɞs��|�t��7k��b_ ψt2�B��p���?u)"WWEB(olkGq����c�$����Q�Tf�e�NE?� Wp5<��%Ұ"�j���/����!�¡@�=�_�h�H����4����\�-s��j�@Ҫ�5��B_��+���_�c���m����,Ob����xy0��Uk��8	�V��sb�L�ڙ�����ۑ�\�a�y�ZSe�5ov�u$�A��
��蝋,�f_J`J�J�4s�����TO��N�w�ɖGUŇ+KF�&;�Q	s���{*[K� P�� \�?��G�{JR�H	$";3��b��`p�(�]iv��ТA�4�~0�NC��r5]���Yt��K$��Ɵo
K�q����RK�+�E(���oi�q�����������'��q���=����7�u&ެdw,ɛ5��1���Lh��@ �wu* >�"X��8+(���TZ#�a�?�*f� J���v��rhœ�%l���%�Ź���T7_y0M���X9��
|[��JM�f�Ҍ��E�ޟ���!X�U|}��'�N\��2��>p�[_��;�{�	+ޘ^2�9��R�k���h$��j�3R!� �Z��V4e��'K�á�Z�w����-�2��e�8�~�\ͣK�3R�6���o93׈eTG1g��t̰��!��+=��j:���}��ӵ�N=o�H�(�M�3�d��`x�C�|;T� �/�31B�_�|�!���2>���`��R=�B���6V�� ��d��v���EðR��������֌��ב�п7��P�47�
Q������7���5d�;�ʽ��f"�.C	J(yj���c!s�BX�r�����	�w|�)�&�P�s��c�fJ"���[ɋ�6�]��_��,Ʉ�w�	c����������Z�x���LCS��j<KTc�qd���&�m���iJE�J��;9�;�z�����MLFh ������z���|`e߮ ��)뼉�;�D>�y�=>)<�յ]j�` l���eS��k�	o��0���G]�Ԩ�����Ǩ���"��_��_�m%˒��N�$v�k��4����vA���ydҥ�d�����*xz��vA�]�7r�FOy���d+���S�8�.�{����#�;�op����?D�5�[����S��Gc`Spl�\#�Fz��J6 t�u�9�����$��R��:�K���%�`]�+���Sf6�Cw�?��x9xD�S�?�&�h���,C|`�&�������s�.�t� 6�(�H�{,���hΈ`���y)��wb���Cǰ���A�dCWy�f
t�"~?��T�б�EU�< ����P���3�śڜ���a��ٲPA1�(mBC�#�D������jn��&FXN͉K�S��֟m�5͘�wC�q>vl{,�Uu��I�s֜�-{�qڮ������6�$��{́�aށ��(�V��UZJK���/�k���F
H�d5PU]�@Z�Q��HP� h]�H���5����:)�!%'h�g;v�A�UT��'�ѣv�h�$ �F��G�)[ݘ#�._�� ˝2�J>H�KG�D�l�"R�?����n�e��ӟop�0g [�f�}���b�?Le���S+�9�4��M��5"����Qˤ�M���EȜ{��Ԝ��{���T-�od_�Xs�6�	LJqf
�k�d՘���Z/�xpX��@���\C�i��jY�:5��&O� �o���� ��bO7�XJ� w>���z>�2u��t��o��50ï3�Rv+3�`�"u� �UD�I������rO<aD8FHv\��غyHbq
����k�\0�NM X���I��~o�}�bq�Փʌ�!@.\nT�����͝_��dz���~G�L��x �U�M#V?��nS���_�'Z %"�:/+�����֛��j�y�5��HTә�����%5���_W���a��χ|m~���!!V;�/�d���b���(~أˁ]��Q��c�2���.}�Ԡ84iOC��7ߴ�I1tc\�E��B9C�Y��mm9d�b�.�dʪ��J�j�v�N��B�Ϥؑ[=�򗱯��Z�-JG~v^�C�����{R��l�y��E#g��x�M�}(5+J��b&���bĹ{mV��=�xo�@��E�,Y�2f"4yn��BZ-�Ѫ��I�X��5���F�����O`��џ�Iϵ!p����Mz�s��A^�2����qf�y����S#������)3�.��#ޜF�H)��轊����:/���7UN����f��\�+�Q������7���bN9K	��

]�⯤e~�p�cym�.Q=������M�X�\�}.��1�6��|�CE�N}0�ͻtDt1����I�]���m-9J�&H�K-8�ڹP��>T�H'��D^�Ux�gd}����C[�^���^�0�R�i�s��,{E��:캷�f������@�-�ܧ�$�H�D�����x�=c���Ay_�M�<_
8�:�
�%]�2*XD��w���i�>���`p�$�|)W����W��� !�\�Z�g�T`4�t�P�E�R�8u��x~%�d&;�:7�u�x��%���Â��g_�Z:���Q��Ӛ9{�_+���̽�f�u�U��?�iS��zA�Ԝ5�	&Oӿ��鄝��3��f��R#�r�UF���T�8�a-�,���ϖ�����GuT5��L�	~w����	x�Kw���M�E����ZY�'dn4�Kǿ����dst]��ː��$ �8����LO��ʳ S����,����q<����c�?�3�t,�<a�Y�\I�d�d���s� [쿉;�Jd4�#��[kŢ���@ ?��O4����Ѫ]��8�$��V0���ߎ��s��ʩ�,���"}Z���ݢ�n"7:���n �:zh���ތx�?����Y��~�X֗^?�?aq�g� ?��A���u^�f��x ��t�W��_z�0-������6�"�f�����K�h����{e´t�h�zg���f�1�@&q �Y�)��I��^e���U�e9D����֙~,��^�`��R�y���~���	)�.;�n-���.s'�gs���|}�c�z	�LuY�����񯧃k��seo�:��	КD2c-����)6���i�	~�O<��.Q��]���Iz/����mR�{]�(���ҳ��D��ٗ��w�;4��d���܆�@KÔ��g�ƅ�p�rᗧoڻb�L��ՠS��d
Lj����7Յ�	�"S��s�|��#���{N�%��sPOp�s���,Vb�= ����u�ۤs�!�Ռ�ɖy�)�C�Ƽ��\�����]���L�<O��1���X��=�)H��Ƿ���@F�G�?l�Cx)2[�����$+!vk��^H��'��ty��㐄�d(ܷ�۴���ҡ3G�d�:�m�L�ồ�+gRL�UD���Ȼ� b���"5��#I�ڜ�t�cr����$c����N���p��"��o�,�.z�#ÿw�L*#��sm�����g �Z]oq}��ڈ? ���Zv;����DT�9��B��S
�+�(�0.J��H"��5��y�\�j�O��k�n��#�^Q�Y�rǢ�R]���3��Bn�5 F��r���d,/9�-�y�����Qh�R�Гv���y���o�B��)�I¹US���+v!��]���z3��
�/�9��11���X����7�k�u`ƽފ��↋I���+2!s���;o�/BP��ى��>�{
`ֱ	㉸�0�~z�Y��(�! ��.^M� 4�+�sj���Ԅ��{}�:N%3]Q�3��|�@�Ɇ�<InPr��[}�Vo�%I|fo#��UhpL����
.]-�7�~��{�{� �Fd���ݔ��sod}5إ���+�4eQע��I��<�|��!���V��ڤ^e�)�gb�Y��L~�6/�*��3�3��&Lr.n��VD��v�[����#��4���6J�%����3шl!!����{}�����͐k�;���_�a�/b�ꠐ��O�f ��8_�R�+��#�8�����>�p�O��pv��s��6�F����3��@zM"JN����i�}� >-J�b�4��;Nq���K���(��i�&��W2���7φ�������K(�at]�0������U͈�]�ۦ�-�VnWj��\H��#��ůM$�W�,���]1��S��+�Q�DB�%J�ݣ��f'��,*��إ���Nh�׽�GK�w'��{�XO&��+��Ұ �?�N=,(�~�l�d�y����8�SQ��8�nw o:o�n�h���lB���{��@��?����jAyX0����f���T�Q�����Zv$[����$ --A4��&�� p��5��n��ܔ�L�;H'27����sȭ��@<��>V8�������a�=�C���0�Z��=x�Ջ�6l2���W�ã՝@��b�z������7��v�/�#��rz�<���1���^��8��ѿ��R�)$t
d?���^r!�4��5#����M볢4��޼-��s����Ӭ�LB!��g�S���_�C-��^�2t�����z7�������r�- p��<�X#�^���Y�&�joȐ`:Gb��}� �V�of_ܩ�I{
F���p��N�4;#~g�U�^��IqsB��1�tILQ�S������o8�y.`��7 �o�0��'�I|zYג�,�B�����Nכ�AZ)�\9kK�&"�ST!°��P1M&��P�8c���6�PX�=U{x(�u�*����!$�G�Gt�f ����P����p��+aXTD�fƻ�|��0uW���f��!����M���\,�$]��@�'�0�)QF
�pυ87*ؠ�1��p
���� ݖ�/�V�m�e�c�*e�;5v��n,��`~��"�y��S�rU��S��v��	f�*�1��$'졇��'�S�q�U���uo�7���;��g#hпnV߅-��f.�c��'�"�S�m n�_�yk�˷�V�W�Ut��JnM<��U�s��� ��J֖JLS�,��02)8�`uph�k?%}e��1Zƹ�e���k{�s�[=6V��ǳDRrJ�env�e<0X��S#SW0�
���)+�a_)d$2����Z[!�S���!+��0_�2��&���#�<��,�m�+�y�p��!b#Z���"�����kPx��rr�p�5j��a�`Eo�a?���1���o2����^�/�=�Ծ��&aƦ�4L�I&�W����9�%wLt2|��#�~+��7&h��_ع��C�-%�ȴd��>Sh���Yb���E��:�ǎ+l�|g;E
�P3��nx���⼯k�=�J�7psu�Y���.0Ed�c`�>�$J]B���iQ��ylg��(�86|�|�YGQ6�C&_!�� �3��غ��w����#5k��R
U�A���We�'���.
�I����U��ݴ��2-D?�-=���c�x�ġa<�}f�hO��?��+Ef/�	�eRp�����G����={7r ~-{�0}�̿�l��)7i9���s~O���/��ѱۅ+��#�>rb{t**��T7�F�ma�-��d�ٕJ�h1�>�e��_�dy��C�Fr.�b�(V���7�ҍNR7  �T�!j�'�����6����ȐVV���D����_�����%|�z���)���J䀠J����ˆ��U���}e�����n�.ET�~�g�҉�8L���%�E�5� �DC��	��֜&�
��ԇ7ζجE-#?����t�`��h�0��;Z{��nx�;Md#v�yO��Z�<�����(��s҆вk���/0f
�'/�)(�ە�w�6yHe�W-�T��/L_x+#B�T�?L�lSW�amu�#�ɂ^ ����{�`�_�]1J�4:"'���g����0_��ME�j���J��l<��W��� 37�R���L���%G^J]�p����B��Ʌ>��(4�����*T��G^U������u��K*�S�	.*Bd�=G!�ϓ��[��l)��l��V4�f��*�	X�s������o��9���G[��qK�U���})�Ƕ`UOb�"��/&n1P���}�6�r٭�.�n�^x�|�A	x�"z��Z��ӗ���m���B�����(��b�E�+=Q�XҨT||���*�0G�|{���n*�KGQ������g�V�;r�hNM �l�;릓��\>�o�Z>2"��'��!��$�9�A.�S|X��Zr(Rw�eL�ꀁA�$�2��1���@ڀS���p�0��^�����{ޥ,镰�F;�_K��(rMp�UM�Ѭ e`/'����*���.���q��<�mw������Z\�DJ��ݓ����؃Q��jnI`�x�}�ۅf<�e�y���ӍSe�2t<5�<�z'�J M.���og�vNu �@Z����Ļ{��`�:��T�?��mOV��$���P�å�;v��S0����ܼ:���E�i �ZlG]�=%�卾�V���6ׁ:!���V�(��*���������kۆi���}�YSY��#�����i�_��ʈ��5�<�-��ي�	�p��7X	$\í("����z�q�3oA^�D���T����o�����k�Ӫ� �0�[����a�X��1Bh�������j�
�-�t��<-tkdT�!��%��a���F���O���&�}Ǌ�������%PU���$oѓ�ԣ�����ߴ�_�-ؙ@�CF�6aЪl�{\�7T@1��e�!r/�悙Ѷg���2	MV��q��"��+�FE���gv�Kp��Į�n̻�=؜��Ac�u2+g�ؙθ�{��C©�x��_��cW�.�$�x�2�����/��且� ���9:��,�E�U�C�-�O ��a�.(�����!�Qz�A#tUc!qʌ��d�+�8��{E�+��J�:�>l$Q���ܾ����9�,�9���#j( 9�6� �u���&�PLO���7G5��Ls�I,�p#�G��V8A��i���Pn��t��~�WI��(jbj�i�o��HR���P#��|VF��%w1�\q>_ӄD�U�5
.�E����~�~W�G5���R{�E|e�2�L��YnF�8�[�ήk-�Z������nf��д��-(������ڄ`1��-ςWm���F�m������L��tyd7֨p�����L����CT�|l�(N~�X�R�w5V�E�z�]����'�5�Ld+�5X\���s&_9W!S}_�VR�`w���ۥG$�n��]MC�ѝARB�����8e��7�:�NQ�������H(��9|����4l�k{����zH뒃S�_�y�����0�g֭�SjE�>���z��4��X[���( ���v�6Qi{p'�+?^�0�jD�{3�Q���_Ut�50g��q�W"�V� ��I,�k�Y���ɲk���L�)f�g6/�X EY�\w۠��V,#q�o�i<	�6N����D:,)��J�b � ���@+��=Am�볍^�� �ܭS|�EGs�W61����j��#a�U���7%6������gY�k�1`5����rmd���Yu�cQ���[�:�)a�z}K��<��*`�,GdtBIPK"x���շ�w ~;�q55m��bY��7D�a�N�e3��X���K�?*�?�
np�F�J@ѥ���]�H4� �t�Y��A���LA�Ӹ�Y�\��a��2c�r�p��o��5E���Г���{�T	m��[t��6y���A�6���̂|�p $?����5K,����jZ�>Sm�ΰ�ht��P�JVZG��%�G����2ʋ	�y� D#]��0�AJTL�Pǿ��1��8����F��	q���[\�]_M��xhc'N�����Өth%��-Ll.�t��޻�{������v�K��?�]�e��ή��@̩���P6�㭑�S���e���:}��2$��.c���(P~�xc��Ҳ�n�"�M��Zmp�{�F�E��(�
x��ľ��1����`b���iO��]H��?S����-��'��}����H�]�����@����Ή�+Uc�Q>�2/O��k,6�������m�9@$>��?+BD����c1���ӊx�SSSՋ +(�?Ss'�5Q�8�����ē�g<2�U� ��M)�zPB��M� �W�-���3�#��(����� 6���$�$� �bb�jv�S�6슉��	����}5�1HZU%�mD������L�V2�A��XTo`�HJ�����wmg��K�w�H��WѴ�.��F;"�����'\���g<#��~}��]�pi+;J7_��~�����j	.�:#Ϥ�iOz@���I�Z��dFcÞ�go<m[�xջ,_&�a~$F����$z����g�o��k$k��/1�
r�ү��t7�*��2�9�Q4}�A���g�D�۰�{��$ Ss6O�Dp����A\V8S��`^�Z�Q����gW��|�C�?��xF��Qi��	NSeo����e����ܧ���N��de��\�(�I�ȥ@OK�_3����+�� v�n!���4/����"�xH�U�L��*]�<N΃�Mጓ�Gw�ne��
���{;�������83��A݆3H�|�����+�l.�
����n����i"��KE�y��N�~:~v�s�/	���!n����g��a�^�/j�7y�z��H�~�<DgJ`��|��x\�S�g��;�u^��_Yؑ����;�a2'��쌊�P�����>�f�(�[�x��$��T�����"mn��[`O�*q��&7
���F���:�����	�m�UA#�6���zu]uU:FHԯ�!�D���A�iJ(�.�^+��Ii��dfi����O��v��6`�H�!b��z�|����|(p�/]����Uf�4'�R
02~����hi�ռB���0;���&4j� 	̟�āyQ\`��O^�����4zI�b�tO�d�0�����r:Uo?������>���A�y� �����¶4�z��ȴ�4,�^�i]�7�^Ӟ�<s��.�@k��h�SMa����j�y�Q}OBt�����<աs_��ȥ����'�y)���g-U:�����:.���]P�4��B2_�b�<���zל.�.�Á畒׆P��� {��5ʊ��f�	A1o�{2ʹ�����"�\�pD?��= ��4=���C��A��LxT��V�
A���QW�y�0賱8��7#cF�E#�'��v,�� ���t�ӣ=^�ƻy^�5\�?�%��{H�ʒ!"�T��Yo7������ؙ���醩��+>
���F��j��-���3��=�0�0ܼf��Aa(�=� ӕ��
� ?^'���pއ�� ��n�[IHn��7��u�w7��-mP�״�G}��w��sM�}�'-�&3�oAH���!g�]���Q��ʐ%�e��	��1��'�Q?J��1?�^�$6��A�c��� #���w� �?I���~��~����2e�EB|��B�b9��<��G&�S���G4���(��(��&�}�$$�����>$p:��p�]��h i�K�ӂ=�p<�����X)��{�[χG���X���u|�h�;��[#��g��6y
�\�v~����@�+��<d�*M�<�P���-T!�	Q������m�˰ۭ���^a
��w���'c�m��ם-!~V{D袀a��Q��>5a�+1"G����tfK��%�жs�_��OY\P��
�~ф��JC��¢��hbT%��h�e�dE�fhu��4����f8\[6)ÿ���f$�	p?fF����[^��Ten�՛� q�4?ʇ2��k�Ҕ"���5[:�u3l�S���J4�?l�k�`���Ĺ"z}��"h�y�T|��(p�l�Ųi��!&O�؝)ht�����%4_Ye���`�uvy��C�I�6�6��ח� ɚI�k��u���[�vo�v8j�t,=��v�0�m�K�� �uٜ����tO��8x�"]3ޑ�n�����"�]�?%��D���_�%��'��)/�L��<O�n�?��ɞ�KS>�� ��@|JJ~��hM��J���]���O�f�&���{����17��5��#{6~1�1��"e���{;VI��q^�WY����h��ً�K��k��[��I��;G��\jS�O����lj��)Z#��$:ӈ��C���"�����T�2=���V_r����)3�8�Q�؀�9fX�����0s�XO���F5�*�~.��L���`/7C���[��X�L�2=��W;Ki�)��ǟ2���V�����iz6�nb�շ��>�A����Ќ��oM���[a������ckKn:�*�����6l��}�.v�cicS1<��aWU�C��L�����w�,�rUa���P���w���/A`���-�=mr~��K2$��Ɠ�{Tp'�����c��V�4���;��/��q%n���JC��oE����'|�I��:�eI��^��:���\��1D�-����'�S��N�{W�� ��ߓ��>�N:-}�f��N��xX <����c�����
�d?�% �vPg�ɯ^z~ö_K��}lQ�E���=5�[���'�0��Y�T�N`ΖM�y;�*�C#DI��j�I�5�p�`�T-�=yc�����e�K7B �ї�N������%4��<'����Zi��2�?�,�~��)ǹ�)�Y��!�p���
i)�+�,�߉�T>\RWVz�"�R��~�:�ʃ�i���k'�a����<�jpeY�ɴ�l'4\��؉���CE��m��I��8��R)�ls�B���PI5�,����SA�JJ*%.�R���0ɿŨ�J����tA�0�1а���ɶv�F��v0�H�����+�gm��I)�U2t�;�Г��MX8�y�&�w��������S�\
�t�Q��MQ�:6CǕ@���&�9:�Ny>k\��;i3x_0�1i��u��*��7���>����&Cʜ�p���d��{����v��!����c�y�����z�-Tǖ�_�'?��|��f��m���yh��ˡ;bܶP�AK��i5|��0�eI^;��Qy������J�N�����o&����X�T�I�Յ��a��͟��(_J'or|�ȫ�jB)��U&l�q��H��n���Yi,�M��Enk��]ѣ����G\}Rc�FK���8�4b]$������������`�w47��u�pl#���J�SlHUn�K�mP.^u����,������yX��ќ�4�d���eyY+!��>��_�Ǧ Q0���_�������Ur�g��w�$��d�f����	x��F�ϧ���Nq
�߂���,�{L�v�W�,��/LDs��Md�XML\���o��/*"�N���r<�ˎcL���{G>���|�������̌W�ӫl�d�l�^�y")+EL���$�bQU.L��m���+J�������׾?�Eq��v��Eo�Rg�hAԝ_�t��q���EVpZ��u�������>����JW���8���0u��i|M�P��
.�CWB��	"���t���k�c��wyn�_
x��.��ɫ��� �jġ�����Ё �Y�{�N7g�t�\H��<� �+m�v()F�ܳ%��,��}��U�1(�O�r�_��~�7nt�R�Mz��E1�"I�o�)��|$}I��x
{M���^c-����fG��!;fƸ[�(�ۤgJd���!�&�t�>��7��t!$;�E3×�)�1�Hh�`�u'�6r��j���B>Ȉ����y����Y���QX�1��,�W�Z7�4���N,��I'�ur��Xi���+<A	�_����lA���6=�L9zz��j�"��o����ղp�l(��T�"G	X ��d�Z��I�|4�w�8v+X>B@���d�	�ݼ�Qq���q[q?--�%���]�uZ�:M���e��k�z�r��wQw0�`6n�#´��o%w#�'�����wL���9�-�����;Ժ���ﰑ��+� 5�7RH�a���o:�e4�Lȷ�2��/��1��<I9���)Rb����}Ey��(�x�2�Z�	�9G �L/��3�U�3Ҍ'�}�UJw�BF�:���zB�%.u&�����ѯ��k"�M�C����&K����wvEa�y��/��B��ѥm�,w{|it�L�:�~�x����l��J�����f��EJ�+�sG��'�r�����L�#��n�2��]tq�� �:��|2��'���Ah{@](��IŜ 	b���X'M��
�����:D�JK̤���?��Z߿O�̀�y��"$>B�Tp�<4뀢�oֵD7a\�Ŏ��㯓1�չ	ף��y�S���91D{�=8
d�2���ˁ�[�ŋ�%i~פ���e*W�J�M��'�&�h2.�X����2=.r(�W�a�X��R����B���� �a�5?h:�TU��̈́����=sp�~ЍB��HQ�4s���lM/�6�69�IC���+�����L���)sn���Hs��s)#�4���6�6��'��+=�KOkO�{m�3��\=B������}�Ơ�Ā�:�J�5�="��ՊS��-X��������m���l�o� ��\oF���-fW�i>VfgQQ�;�cM��
:�<�|�����7˰"G_�j<����}��orP����gM.;eIu��%�}��tJ�@S�����V��/=F/�
�B�2�E��@[�O���[�C����!�_F�q�AhJ@��f X��؀g�k,�~]������wF�a@�c�O�/ Om�6�ݍ�%��T������Z�����E���Յ�1�������Js�pŧ�oS.G%��؆m#dMU�SlZ��MK���3_����Әߟ��K`�{ً��,M�J0�[��O܁�����g�^�rJUG���f�:�,�G^6�\��>j4.����W�%�����`�����Ɯ����?��Ө�}��L�t�m�>����|mp�������I��%�r���=G�P�=m<�����{`-��:S I¨_�~�X���T������#p��	Ru�{��$Q��×v���b.>�2�6N7�DP|	b\�$�b/6e����k�x�p�
,1vIk:!�C�k��n�&��II�h_g�����d���/���x��5�ʪL�xx���6$d��O��Άj)R��N���I?r�n�d�K���,������X82DPB��e������_���5�١�J;�B��|���y��Ș����EߚՎ�!�`��l	��$^$}Hx���nu]�~Ck>Z@�gJe.�~��s}��o���qm-,�Nـ�z����
o��Y��*c@�B�b��?�3��	�1"!���ɫ�g�?�Ta���!Ի�J���D�Ǽ��tM@15�λd}Mo�M���S,������%���#���ֹ���-�� ���ı�#�F�K�u l�y�(h�n�³~A�w�9%�����sRQ����&���k�X?�;I%�&X9M,މG����T�,�4�h�S;y*�j
������<(�p�U0��ҥ�$4�Z������������9����|g�Rl�y�����@��ۈx~&B���+8ne�p�\lI���N��~Ӎ�CS��J��ߴ�v(W��{����\v��	]��+��m*����ѻ�>�A�^�JN~��'�( z��>�0��������P�8���J�E�11,q��l�s�#��a�3�O4�r|�2`�JI�G1-%�i�mǍK����>"	�P�U.`��@�z��d��*W�~1Ħ'NWE��;�#'�1��d�#Z:�^�q�9
�K�[f�JD����5�ʁ s����at�� %q,I�%����
6,�'�m�`R�?dk�|l+⃟ؾ*5&�or`3>O��DM�h�zoM��Zi27I���f�t~8��`jmA�M�WTH�k8�K����8��g� 4��ۧn���������T����Fe !�e�s���VW��FF�u������m��Ku��D%�ep��Ff�z�b�.P&�3폿̺8��!�p���j`u�Q�[�K�}��М����@�|�u�
��)��@fWI�����:�N(����H&�L]Ɯ[Z�A"]�U���I
��a&���η��M.q7xQo�ÁGY�f���/�oH6�EEc9�T
:��Q����ΔB�ɢC0%��b�+���0/�q���|���U*�v��wl֟�J�/�e
l��?�O��6:
��,��QO��ă��J�ZH��K��Qi�F���]感'�ǵ0��Z����t"��1���� �JD3��lR��K�㑵�h�4U%�J)����P!�l�^0�rT��Ӳ��1_���;VAu����'�ևE�t]
�cƩ0uզG}Y��U���y^+�D��B >�b���9��⛇�T�e%���a��7: �Z��#Ԧ=��{�=l��pP0H�U�b��25V['�����1~�� vIDZ:a �0 ��3�A#g�#rLؑ���N.k���G��� ��fve���d�/�9�r"b�y&x~���M����(�O����O���o>$F�j�C\U褓�Q��%�XSiu0Q���y����h�z�M�"�^E��LF���*睁Ǫ���DFH<i�w�ơH�Z�s��������qxj17��a3���6H�S��Ŗ��U����}G�G`��;+�K?lK��g���ɵzH�hgEɈ��"J$���ڼ�IUPjho��G>��K�V��'l����'s�*).�Md�ty_�7x� 0DK��q�=���� 5�~'��:���Al���j_]C� 7�q�ā����+`����3s��7��)����"���G�џ^���.��^!�.�[p��O�+Rx�P[�ǿ���ѠF�(
��E逯]�P�aL��H��4C�!�Xl�~�W�XC��ǈ�5*��A�i��J[X���3!
X]!��^�HG�"���갊^-�J �Q�����*��vV��x�#�<��ܽ�>׃�F���D2���7qۨ5�b �P��E�>M��� +sW���oh����+�%6{d�YN��Aَ��|�啭?��]�o���X���_���)�5o�M=��	tڿM��m��SBA�׏mtY0�(��W����j~{����  �h�a��+R��b�j:�L�'�`KD�q�=\��E�o.6G����7<�H�x����WH�Bql~�hUWӅ���y�h����v&��A-T���~Df�'%g�?`X�v��G�mq�r��!���,5�������4w��Ј��5a���J���	@��e��ͺ��N�����]Eh�;�/`��k	��S(������y(_0BTl_���H[���%_LrY�j՞���c]�����nI��3����<mq��7���m��!���1��L��Mc�I_�� %.cޛ��3�J�y	��s�2���¼�L�Ļl��Y&�}� R(@�y�3À���H7��{,�9Jo��*F ��>~3�!,��Lp2\%�_#�=q��ə����7i/	|�aB(��Li�mf5������pđ��m�"z�9Y��� ����{O�0�$y)�B�d�w����'�r�����"���M� ~TN�l{K�a��*�'&r\��=~ ���p�}����|��/�%�E[�����;ul�B�Α�����l��?��7��$Pv�|���T��'(ͣ�E��F�,��5�:%�d��H��}	�(&����Ƶ�ҝ���=K"�u���6����9"+@"�������`�Ae�,�&P�C�K��VӵD���C���r�6pa�;�����!�E��=�[��qsZ�Ǳg�I%�>������D]��;�5
HF����ψN�<P 1�0f�p�$�V�GX��*r8V�L4�1/]�G�p��ī㺞k��ϋT������O�%���$ƥ�`X���-�haO�~.��G�NY�h�����7�Fa��0@�
*e�H������+e���"�s7����� {��'�q�~c3�ID��^��X4Ȉ �k{}R�4�`@��Ф�X�N�5��>�*��]� �y\�N�8�^���0��Mj��c�v�e�'�4X�,X�Vj!)�_�@.(�������t��2��.�7��%�b>V�^�/�p�*�`���i-q;�i�>�Am߹k�L�~�?�p�"���G?����u��i���6�ow���ؠ�#9���^[��u����Z]����!,I���4��Ͳ׺=�;�6�)2�
�D�M���G��E�}���.|푂WI�\�6A~{ׂ�n��]E��U_��~����|~'�I��j�ƢQ<��>��C�o�Q_,cG�-�a�xfΰv�P�=�A����-=5c=�PW�W�/؈IXz,EI��5��Ƿ�A����Ъ6'��]o g��1�R��*{��㲢\Xp�����s8�Ęc�ǭ���|���]�����g̋��vtZWF�Ђ�@��j���$���̧�!�
;��**����ҴCԊ��,�<['S�E�`��;DR�V1�-��)<�	�"��4�Y�"�(	�����X�L�'W�d^/��m%$���=�n�q�{��� ��.o�ͳᎄ-�@�D5��S�T~��s1e�XST��m9r:sӛx0s�����`���Q�ឋ�����e�o`Z�3�6�\�ަ�ȏ'���Ho/� �ސ����������+�b�JA�����i�ж��pc��x����;ڮ�hm�ǡ����B�,�}���߱Ù�4G��^��{XىH��y$���/XCI0m�x��&aTG�+�`u�rv~UC�,���9a}�^�����Cɟh�mm����� s��Xq�H�+7,YR"��W����_ �؇��{ ��P��;Ş}sź̝��*Wkt�Ak�e�����y�Z��a������f�����x��Vٓ�TM/�j�XD+�i�M-��72=���ڻ��g{GSÎ
��ɚЦ�}��S�OX�KL�78ޗ��@.�� �ڍ�pu��o���=D�%`�CH��/� ���-��!���7GkZ�1uԙ��V��ޯ|�F�"7�!NQ��أ�� ���s�8A-�&}����_�BOr�'�~��C�[��e)2�.=��~���s;%��|6�v*�!)E91'Rzi!?1�RJ�J+�� :�/��v�*�U.�S�K	o��A�JL0!n��OA7���DY�q"�و������� /�1��A�\�L~�M@KⵂE���UK�y^�a-�Ί�rb��%��M�=�ygt[���+�����b�����: ���`���o�s#���`�&���Y��0���͡;��#�`�
��2��B��\Æ��]������v~����-��TŴ�y�A���23yI�{��ɞR�Ȋ"U{F/o��;nN���Ͱ�U�s���E��=�H���w*y�jyX�A��5��l��w~,O��K�h�����(Z��$��r'��w���٬�O������,�4��	~(��ڍ2� 5�5�!���;�����Go$~��,��ǉm���e��n�`8�����>����%�3�����8��y�=�\�5�o"�Υ?�y8��ؤ��.��/:�]�S>�'���3}FZ��A���N�f�0����1�6�Yj��l���R�m?�y������Li���ɵ���/���[<<ʚ;���œUW�8�a���:�~EJ��{N��d֘d
�Р���ei�g�����o�Zቈ֥#P�X]d�J�r����P>��Ʋz�x����C��c�!��э�[4RK1�<��=�t�jf�C�2c��K4�2dQ��	H�4��U�,�&$�H��b���}(#Ziz��R������"�k�v����v�plcx���+]��Us��ț��-����%=O˫o���@��F�Fmo¨�M�?~�^��{wfi��,�n�.d$�m��:��2#yS_��&�m�3�/k�`6�Ze��pL�r�*r��A�lx���?��(cRז䬇vҾ�t�z<� �G�F(�lWJ����\I_1��~�'_�B�i�̑��0%�iӳ�wu\�X찅'Z�n��T_7&�X�����t�Y=�u�Ĥ�ُ��� w�aU�o8Be!�-:"�]"�,B��y�d����р?��{��R�ͨͿ��K[��B��
%V?|�I}��y.�13�OOuJ�d�^B�oR�V���b	-����^k���I)��c"����I��y�ɋ8xyq��醑>A��[A���\G�>��Y9��]$
L�I���'�a	�xP��[��m)j�!&�4L��9P��<�T
G�3T3P���<�#�8Fۼ��-L���3]��YAh63��]�LN�������[�����م��S�p+o��Is�����f�PG��1�-��������pagG�n,ڷ.�aG�!&ʐ�c<v�����&ˌM��M�5����=j��`�o&�#�[�';�������0����f#��x�Ɇ�Ҿ��ʠ��¸�i��5+���%��0
��4��`%����l��&xW��Ա( �}cmO�I��^�T�<U�퉝]� �L���F��:D �[ ��m�U?�2����3=~�5т�"E��,&?�����P8ߏm�v�R�ga��0'��n�������;��O�0e=�>� 20O��#�u3<1p�-(E�Yl ����9S�{�����_q����� �Ʋ����q$������O��\<�(i�~%~Ţ� �)ߩpa�h�G�`�Y#ڳ�Ex��9�sݙ��n}�E�W����S�5��Cvy��S�XyL�d��飕�e69�B7o\j����7��{���p��0�>����K�6���k[�Vg&���Lǫ�3�B2#�Ї0�>{D=�wm�� �8����'_�T������vW!�"Ќ����Ä 7X3�|i6��c�e�pzzv5��u%^���9���o�S�m���٣�
,u�GhF��!N��� ��=�E���J�Ӽ�q~U�2u�X�4�\�9�{�<l�����?�i���2��.1��+/p�\ ��j�;&��u��W���-ŏ��,�uᤧە	�RxT�;4P!���(��2��� �PgߋБg�QuΣgEw�>�0;d����υ��5�=!�͓�B�k	����]�ݴӚ��փ=��X�4�,��<��ft��eQ�f@���t���$����J�o�CiyQK[�R�!A}�g�$�V�#1樍 {�V��S*@��蠯�C��!�D�n��1K�"�±[݊	^���s�N�7�ہ�W�Y��N#HG����O�#Ʊ =ڷvRWi�,L�^�-E y���A���њ<�X0��.v�b�~��o��FE!̯~G�;ۡ�hH����K�ы�S�L�H����@kP�E���'��ڽH��SH�W��pI��頠��R�r��}���:U=�㗆�|x?�ͥ�老s�J���S07V��@�͛#U���R�7�����xV��.��)}���}��do�@R=��V%Ԟk���OB�ޭ��B��
��ӌ�4ˣ�/��<>��Ǧ��W���$��ü�Ii)�x��D`[���Gܜ
���� �2T�d	�
��]X>=�t�9��oʪ^O��]�N��X�����X�{	3��̽m)����s�  ��/��o��!��զ�M��7����[��8�&�P���u�Zia���&.DR��θR`�rŠ~�i������&��"��Ɂ����h9Skհ�BJ�m�E��I13�K�P�ׁ4%�UG3��׼��Ei�K[���LB�0o�Q轕�����<����,/nL�V}�2�r�G���h��x���	��l#�t.�T	�H�09���
ݭ�-� Zq,1��������Út�&1 џkBm�5���xD|�L&[Fe�f����eX�s�W���-�M.+��/�9�~������aFXfx��Z��{��1�
�d~���%�|�GEZ�߷-nd>��|`�Iv�{+��FgJbF�`?r�����ȄL��ϠN�n.����V�h*�>�u����3�_,Ј��u���f��Eg�]�B�A����ܻ��+�)T�����������8�qom^���4W���c�^O%JŰDw܀������%�.Y��3Ϲ�s�� �I��yB]ft"�ˇ ��e���_b�]|�	ZL��:���/P���Y��p SXV��Zc����&��߄�R�>{��P����ެ�,~K�V��
��;k��q3N�}3����MG��8ɱ��q�1~5b�nZ�J߽*S]V
+�AO( &n��jn�y�ԡC�ǎ�WU/��-�E.}p0Hv	v��B��H��;bShbӔp`���'�d98z��6e������ �?s/��1c��ك�`�\�����Ԭ�� ᵁ���\~��Ӑ��ċX�`v�0����.S	��sY_o6T�N�X�?�������bV���|��D_�\�b�>#���fzTp�6��Z�vf��!�.��PY�ف�a������w.��"��dT2��Z��#Yo��\�?��V�r���M~�P�#��L�&��q�6"\.�=�� ��f�ȳ���\ƨ}P�he.?뵿����2z�^���[��工4iV�"��3�ٿ��N# �%�JG��ͽi8K�z޳$&�rS�b�aD���I�;�b�S2$H�wW�^�:���z$�'X�AǠߣ�7������މ�-r��<W �;Q6��k�IL��
V����[�"-帅���
]�i��T獭�Qi�9[B�à#�撶��_��|Ӂ��nU�S�}T��9!4Jՠ5�o�J���pz���܆��Μ"�����k��ӆUy(:��o�����ӥX��{�4�7��������
�K�*��U�d\�۬R�4���J������v}�z/i��5�/��iB��dc�V;�%�U�G�S��9��7/��^cI�-ZG]2J�{޿�{��3��u���"$�7�Q(�h�wECܞ�e},Uov�R��{���m�\����4�+*""�>.)����OC���Bo-��i,3��={��Y2<s�"!�t��N���"�yt�1�O�/�j�*��>��3e�T�YC~"F�u=�=���.g�pD����G��]�Z�{@��$��3������t������/}�W_�������UJ�C�h�V���˞���[��p����V�j��iZ�~~G��{�Qo �$�ʲ▸����md��K!�i�h_L�_�r�D����T��0FzD����4��9�Cs�!�5oHl��G��+ �`t���$w�Lȋ�����!ڿsdp��S�ir;/��,��L���4����S�埏 W�W�O�R��Ko �y�Qs�c$����6zD¤gj�e��{WM�ذX��iD�L{ƍ�Ŋ�K��Z|iF����y�����( �rVS�U��6�����j��;��Ш�u����n],Z��N������WO�'u��}�9����$բ�Y��JB��^�t
PX�"��ʏ�v!��T�qk�S��7�u.0�WG�����Kc|���<�d�a��3�������ZEO�M>i���͆�������jM�ל��;��:��\E>�2^7E�j�<��An�\m� �d�r�u?�������}I�X�"j[
%���2}��\ό�|A%Ǝw2���&~qn�T��oY��R�h��D����{�3v����͕�IgGa?Q��x���&A�Ml�	��DQ�X��R\߁u�ݸ�-S�F�X������(^��Q�j?Ũv��/=�g��,���3:��Ȓ����>�Jan"C*�S�	#��#�����@����\�C��p� /��Rx���
�W�%8cz+D�=n��ͭ�%�[�2:��Ku��-�ʔҷF�b|���k`E����ⷪ�*��
 4�㈊g�-:�5�)�N�T�l}���qB얦�栿��
�5Wе�)�ݤ������fq� ��)�_���i]��Z���j$�|�M֏�el��+�Q��B=��	Z���8O����,=xCVW2|�����?�Y<�&fQ�l.���2��,�yVTv�z���VNg+��<��?����:O���4WL�x'
�෈���i�P,�.t����0�}/UHη$��
<�}e���w-2�g�	s�7��$���iNۊ�7� ���Q���Oϰ�HaË��и����������n���	w��.��D6�X�)� ��xq�h=)�*ZM�6��n�4�~R¡�o,�
��p�1y���1'�^R{�s�R9��ɉ�8Yۘ����s[(&��Dk#TM��7x(ݞM盋+KvM��=F
1����'�!���E��qFO�@)��mw�Qf*s_���B����M��,�tl1�`����M|6�w4²�AYysr�o� C'�9T'f$�����!����-H�8kZ.}Q�݀��y���}���+��Y��H������Cκ��
 ��qo2��]_p�������+��Yd�MiQ��8ǵB�ɺ�n�.�[>�������(������Sx�������%9��)�[��~�÷Ȑ�.�s� ��*�R�nz����!��(/y�{��7"���ѕ���i����1E 7h��d�(�?��큃�Ny݃K�v�P��\�/+9��@
���`���OzH�)ʃq�i/ �u{�Ғ�����1�nf�ٶ-���C���~�d�w��8���|�]�Ƽ}i����UcA�d��8z�0�;hſ�춨��h�}8w���*�H�a$����"hN�͒�9S��ɢ�����f��� �'R;�I���."z��煑|$�G�u��'%�ۨƓ|�h����Yޔ\�Y�3�!����f٭V�ƌ�ğ�q}��C�i�F��}��c�#ص�\>%�n_� ~@�we���,����zW�^��T{�z0.�������I��m��rp����bn���Ƕ���ܝXW��f��b��^����n�-����{D�Zo��|����ʆY���H��6��y�ڼ��>����>�&��/��$����͞��wy� �m���tA��@f�7o��v�Ĥ�ߩ�Pp` *c��Q���W#&m��\��f"Eܦ�Y�
�\;�	C꺦�D��˨������˝��%,������=l.:nNv�@TIq�5~u��'�*Z��x���)��?�(����*�K�Y��z�ÿ7"�PF�4q�I��h8�k��̯����E�<�2~���]��f��4:���D��3���K��~]�d�?�qԛd���y+�8g��d�k��ZfZ�Q����բ��[G�1ɲ�ҢZW�.4���j����@�l�]�z�L�b�ɦ�K��W]�3�N8�+��سeU�h�I�a���U�Nf�@)?hy}�*n�h���|3�kt�4��}��_�$N���۟��!���8���<7��ח3�����bV�Y�w�BP��N�uџ��΄���V^��&�y���� !�?O�X�nt	�<{���A�\�	E'��Q7��m� n��_���7���=���=�p�[d�ڐ�ӚoS��rH�א��}�=V�iNOצ���#�A�A�a`9
�#�p�}�g��]�_8~)�u��V>���9���~{Ҽ=�[X5�4K}6�4ygY0P��-�l�� ������ lAS�'�p��ߺ�vpP�>�A,5����>@�L�by�bG��;��]ۣP~�W>�1��/�1LC�K��%b��?��vm?��$sbY��c�����B��3�M��r����X&���w�m���X���I��)� � �zZV��W��@�Q��n.�Њ�q�vd�E�5\�/b/"ƭ�>}@k ƻa�S4v�RB�Krq���@�b�Z'+!��r�iU��k�lL���GS�ZS��e����ڜTܺDX,��6/��m��~<���o���'q�*z�ތ5���ߛ�+mhj�{���	�j��zN�]��>F���5KZ���;<��G�lnZ��pkY��V��e}�Q�e�yݶ��/*+��P������f�F�ڵ$籭
{H8����Z���8�����~d�w"�����M�u���9�\�t9� 0
t���Eof��7/��bj��h+���Wvl;�[����H����jtoD��P��L�M�r���j�[��yn���-Xq�[�k�$��rU��&	]��7�r���N���>�d��U�Fdq=M�ףi�V�/��K pE�d_,�SJ�}r��o�S�%���#.7({93����z�C@�}<�W_Fo�(�_T�rl���]<{�r��ʸ;��@�h�� �/��sil˖v���3\�4㭟�!�
va�k>I�+�`.
���Y�����Dihtw���1�B{���+x:�GtϜ���4\��A����6�0�>�ӯ�H〘���:S�_p��n�'�����2�k`Ng$�?#z�tM�.`ETN� P�t���D�d��iD�{�};�91�����U(~&��Ӗ���.�3n�%�+��6�Ԅ�ϛ�);s'�T�h�q�E��j�\�]�XD`j+B"s�
G�f�@@ZU�gq��k��%��/q��e+f�BN�m��o�S�)mc��Z���@8��@hϘ���؉#��b�����c��
??��$���ˍ�Ӄ��%�h�凾����1r/�sOR,Afjȁ�����*0>��\���
���)H�u3�fpδ1�o�Fj�~.���u)g�譾>�VH���KQ�%w�֦�8�ݚ�����Ӆ���M�����K�9,%�Q9��:|��'q���ڦnx!���;Y#��R���0![mm<�t�̖�(��#��a��0��t�͡񑺪������Gvx���䟏&@yOs��13r�Rm�3y�@�!P�P�~�6�6�	��蕅w7��W?����N ����(�������n��`��T��+�N҂��O��͍��x�-^;[��C�"鑶��0"�����`p��%J}Q�,	������ۇ$U���
k1����	�ʔ�Ŕ�7ٜ��>��:�R���!u��/���o�`8|��W4���h䭀.�忛h�&I!�N_�9Sh�/]���S�a� ,�h蒀�x��\PN&kw�D�]S�I�D�q�3,4$~�!V�PӞQ����tw��G�,7O��7bs�RH����ړ��aӴʸ�iiZ]�L�����#��B�M���`���uF.�E��J[:kـ������c��YR��6���9
-�|`杧�^��'^@��2�Ϧ�M�5Q�	aL���c=��N��8�&��-m ���쏆9W�x��l}�&u����9z ���[B��H������F��h~�Pȏ�Zԍ�0��\��MM��hG���גTv.�^uOL�*�S2.�ne���Ӓ*�֪��9�|&(�\��<�Z�z��� ª�J�V�� ,NN=֫Nk%9zS��;����R_ �
uZ�lMqt�@�;Fe�K���d{pA���%mYY��ycH�!>|Yj��5/d�s�}����������ue�yi���|$�%��2������B�J���	(�r~=�!��>����2JIq�k�`�ˋ�	���y��- ��3v��&H������hnpȑZQ&o.�6o|����Ǩ|gc�@��:���r�Z����>	Hӵ�<.\��&
�OI:�����78�./`Cqؽ̙��-��f�2[�o�׻����﬷ᢤv�6�6qژ���L�i
�|�e�S��\�G�� @�d���#B=��p�r�Q���#�����#`���oX����Ve\��=��,��B��p��A<	(?T��nش���3U}tP�����߿϶��T�$����f�!�N��>�C�GVt1Kw%��,�#�1���&9��l��hb|�����<��B����d{��0�[t\	3P�k�#�e�FkHH�v,TaI��p	Z�)i�N���a�sb�0�Nzc���:�{�tP�s�8\"��IJ��O��2�k��F� o�%��Z�N�K�m)XV�+��A`+�|��l:����d�?,�#�F(z���$@�K䅽|O��fM=�ۭաq�X��NF�0��u�Α��_�,�������kj22��B�
��!�opF~�1!�Rr?���NI9�&��B�ѐ�t �g� y�l����7Bj='�"	,�%kW��ݻO��gjngꤛ�b�;Q�7����ِHe�Ѽq?�u��4����1���'L!�A�dp����Y�,�'�ǈ��h[�ˈV�eSK�Fv�h���@�س�F����v<s��&$��&������,���3�Zv�k�H�b*���,+$.Y�\!Q�Q*�`aZE��.��Zt�>�Qk�f~5b�*�Fs	���Ax��/��!�۵Ļ��S��?z�B!�������D@���s�]��J�k�Ħ��c0R=*_Ao��D0LF9k�'������%�P��Qk0g��I�Ǌ�|9'�~�۝
!1��_E<Q��2{c»�r gV�ʃ����P_��c�F%��R�|Q�����(O��P��ϛCt+���aٞ#�5��p^H�9Q�H����;1�׎n��[t:7��n9X�G{*Y/���Y6���R
�#�;��7�R�X6JȀ�]^=�YE�-��`Q+s��g����+����4b��5����h��LD��N_�w�eeIC���C;��խ��u�EAc����^�Ǝ��wą�u�U���B�~J>f��u_B'�;����1��PH�
gOb�sh�9}3��"Զ��*�_���� ��d[	:h�I��7N1H�LtY6:�ؿ�����/֫��A�|�E��yQ+��{&��$�'��4����@�E�T�P���N�l�@�����n���}�R�~��L�[z�e��3j#��cs�+Ў/V#�}��(BQo�����:'�(�
�^O�|0��z�Vg���&���zY��B5�4g���<��ng�U��Ҵ}ʃ,���w�NK����}��
K� ���ػ
[$\����e� 7n�k�/D�Ѷ�a��XkG�F�"�Vuho%���s�\�ÛH�������"�0M������A
��Qp��ɤ&�Q5���)&�L+��e����fF�(l�V�c8���iO�8��k=�J�3���T�*���\M��:�ꩍ�j��ُEɯ�{��e}��:_2�������yOρO��}�No��Gt��m�!QgY��j;��@��|�z�z_5��ԥ`rҡ��e=֟-�C�(�B:PS��_�{t��R�����+8\�����ф��XP�^�o�b�ݶGf����Y/ڛ���{�ӓ�M�AsU�����w�a�T���F�]�ҁH;{5��l�&���� ��
|��4?b��yv���7�����rX�}ׂ� ����lanL������å�sޡ��0(cW�����TR��;����y����H_�x�A\ݮ#F�Y�Ύ6�m/ P^D�lL"f�=�s�ʴ��N{��*^��%hu���>ޜ�n�Z��њ3* ܮp�e���.BY���#3�V�<$ �?����iEk��P�P'�8|�43�E�A�����a�3 �S�]1����+�7���e��@Ctv����x��k�bV�ŪUb��+�`��q-��5�=s)!�
l0�!����8ʋ-$B�Y"�	���{w��^�{����[o9RǪ����mi	�큒r!���@�� |�T�{�}�E�P��F�m[�&�H Z����Y#�}�����H'c���2�����nh�l�f���g�>_���"\3�����5�V��b�r��p��"�����J�Z��t�JY
"Td�i�,K���c�G�����w=.�C��S6��o��&���*�E�R�f��-��HS#kYiO,���""`�#ƴ|�{d�]-���,In�U���)�c�mĳ�i��?8�XIA��S۝�|�z�%PrB�"Ԃ�Z��j�R��zb����|�GH�EӼ��?�M��zi��w%&l���*��:��"�LN�[_rx���*wAz�ݦ
������ M�Knw��v��a� 5�0g��mX2'�2��"��x<��	��a��a���g� �����/�6��}:GעwdB��OaT#L��R�v��;�n�e�	��<�$z�.y��8)�\1���5�|�éU:N�Q��o���IP�z��n�5��=�`�R��1 �3=�5��G��I i9����
���tW�<�b�����ժ^�
�pb��|�<ly�z2=��k�1�j&��l<�t�\�+F���e��=F�}v�,��g��p�^��06�G���x/�t�\��&_tU�
��S�]=�$�E����#1aA�6��4)�0:Ӥpf��M]�K�cPN���yĊS�g_��H�n�]-Э�5��s��%�~SfLa����'�˚�XiVd�4G���$*�9~�0���6�q㒨��Fn5#?d�} �V���4��U�+�)�F��U������{�_~au�}�4�'Ѵ�΀�f��&$<�a���I�U�y���]�0;���c �/	9x�������!�l� Ny���s
���v�7H�"މc}* �j�5�@	��R+� �S�
C�MB�]7R��>�u���c]4]��Д}�|Ov�$*�b�C�ڮ�C�Fe�=�������T�Q7�Y_V�`�klZX�R���q���e�)��;=�WM��J=���}"ϲ�������%����3�(��{SǛ�C�qW}���1�zg��4q���Qv\۶��(�>l	2�4}�m��}U�'�S��蚛ّ�1Y�)�?�.fm�a��\�H$��gm1������b9ԗ��{k^EJ�;��>�����(,4g�����I0�:v��F��7��j��^@�s�ns�E��n�w�f���c
��Q�K��*!��99�k�XzLa'�H��y�Zݫp7���g=��#H�'�	eq." �h����\�+G���F�\r�������$��sb� ��^��ױt�G��ԦSB��5ec�y�m����+�Q�h� ���`ik�:�m8i���6Ū��d�W�,C[b5��7�Y����ˈ�C�I/���v�n�;n-c��tbק��{x��B������I��������2�]Ru�/}��&��U-j*��� � �N��U[4��mSy�n?����I��5y(O�<=rk��Q��J���"�{�Y�I��3��
��oԚE�1M�%9p���I��J������l`V��p�����<$�+H]^=C���L�H� �@��g��U<��#��y�e;kdy��8Y�� ����)�c9�R8s;�S��K�ϋ��p��xc�v����������&?�W��xT���dͶB��[�4&K��i�YQʎ�wf�Q�D9п�/"+����	!�aܦv���&�����+�]#2�~Ŵ�,,x�ÝB�\�Fx����%��/���|x�;�BI
�
�U�=�B4��́�B�tUFNB�����x�-4��Uَ��SWr@�sX�������#�Fz�;��,UAr����1�W�=
�e���\i3���@�6R�K��6z'݆v�4I.��(����ɱP��Hd����O9w�^����	U�s��q��2��4�{R����6��˗1d@Ρ�n�VR�a�1v�]��\P����W�|����'+is����N�y�FM��6��c��<S�:�M����a��jx?�3be-��XO���-{~Sp#�7P+����#'5Q �P|�t�ئ���, [�*�rл�Xq>�g�En-!�Vӣ��-ޚ6`�i�bj3"���M<٦�<��)d�'11��K`h0ӟ��c+)Ŏ�Y@�d�/i✊`.j�|6�	��|T�҆krf!���v��$B�u���^�[Υ`K��U��PYa��=��
���q�z���/�$`�w'x�s�PE��|g����WY��^1\T�ʯ��i����L�6J^�N0j�Ž�zs����l�X$.��h���Y��st����NV�=���m�R���9e��,���f��Ƈ������aW��м�G0u�F\�  ]�\8�,HN`���oUs-�.4;���ge�
��<B�nSOR#���]3�^b�':C�6!���#��T�b"zEo���o�@�=^V�P���؛�r��(@g��jG@,�U�/1|�����X�1}fH?�L%�f&����.�ډ�&_6z���[�/nt�c����>�_�2X��/�4[���U��@����G�ܬ>�|ԩ ��5U�2��"Ӯ}X�i�����M�q1���irWx�־؂�)�"��6����l��Ԣ7B�rw,���\�,�p��Ke����N*N���],|��3,C<ׁt���~�/�a��|Π��[yVLӟ�Lp1c_�J�Fc
�-;��u�kd�E!��	%$T�z�ܳ��#б�y��s;����k�9��9�=���5"�_S>�7�ō�KzLNj�-�Տ�R�z��F�}V�@��4�6���@�u�"D��-8��k_7���J4$s>��.v
�٫}�A��<�'��k�@�5$f���~ �H-<r��O�ϟ����$L��U �>���-�!���f�ÊH*��6�i��0��>��dӋ��a����n�������<u�����
�&?j���7/���*������T�rP拀�%�<Jd<�Kz�Y����Jg^I�$�WΖZV�/I�D������F�l589���ʝ2��92r�f�-�"�zz�]�tx��٦�������
=1�^X���1���H$N$��-i$�0�c[����O�7vg��x��͓�4�Rlg>s
�{|Jݿ���t~�]��{,:Y�7?�0YVV��T����������SݗN��UG�xS���RfrnȞ�����a������O�8i�H��� VgUؕ�2���A��no�ulּ�h�eL�������N� ��ʹè�[:ʻFԚ�"?rŞ!N%H����]�-��W�]���b�O���H�n!E�OK��'X_��e���1~��D�Pݐ.�'�Bq��=�.�7���Sd��'v�zQ�`�t�@r�k.���Y�Q�X�a�#�����խ[崔�)�sro���U]�bn�&������2Ug#s�*k�KWv����s�*��o�x3!�@��/�̮l+MQf�o;�=��u8ny�1�2�Y��4]�.5��jT�O�@���QǨq��:j��Dv��uT�	l]w���$,�P5�E3	�-�����=�ǵ�1�k���7*m�������	���W��|��ۏCNW���t���6��),��WB�P��H�l�}i~Fx6]Wm}~�����k�O���8��R1�^�/yM�D��<�d�V��C(H��Zn E %�3g+�,��ŀ`�C*_G,F���-�
Q�L�W�e+�����տ�/e��(O����bY���Y�	�Q]�~�����p��zn��������B삷��:��p6�4��*��bC�8�G���[�c���H;�����ճ/�S���ؑ�wۃ�*��ԋ����a'v!������m�VnQ�ѭt�l���)�S��Kx�6�p}�E���8�k�vhk�2[8�1�ܙ˨AJ߃�3(��|�Ҝ�1Y�|�����������[�+��xΤGP&r��z�O��1 U�\�U�(I�z���kIܧԍ��L���!��f�
���aW�c�,�BU-��.J��x�"�Y����#�E��gD���	�r�E����=TmU�y��Fo�{�g$LnZ�x��{����^PovX��q�bU�k�[4�� ixF��+ �G�_��
 L���;|%fNar6�)|x���W\�� q-)&���S����Utl�l4Q�`�N��F`�8��.\D܈2�g�"�������!���Z�Y�WC�qBLE��f�̲��`��%�dQ#٨��h�w�3���MgV^���|�w�(���v<�u��\��]+ l������O��5d�'9x4q����2�JQ���$��H�"^�iZ��ԽZ�m$�������P6��q�n�l�եe1�VsM�1�;�{3���uM"[�NFk�Y` ������a��d<��y]�T�Û��[ ْ���*f�;6fR�L!�� OG �U߹�	�[��C�]�i@��Y~�P	Ej!4�N����|_���@��/|_�K���WɅ	@b��<��:f��
���چ�kɟ1U�V"4���.�	��=��ܘ���E�w�b��u�fa�	W�NM�hNx'S�o�y���$�J�.enb�_���m�7)���a�ɶ+�"�u���~`1ۋl�+���a<{��K�`�XD����W?oB-\<�=�r^�"zF�+�q�R��:?ui��D��+��_��GT?�5�`��Z�`L���"��rQݛ�:Ӕq�a$�b(��E�갻?c� *k���U�o���������]X��j�1Ǐ�#u6$rN��S�@�{������@�SC��A7Ʊ�"�X��;K����R�6�&\&���ࢵG��28D�#^/��_J޲Y6��I,�b��k��gՀ{q��~^*H� Yp;髊�rݚ�>��������y���.bz"�!U���;Xs^���^���&@�e����0����H��G.m�ȪE�\��)�Z_�A�`���6Ȼ�1�v�Qѫj*�i�jc���LC�h07�A
��&�,�j��f�AWɉ�~���v�ȭ�J�Fh�WM�g�$~o"�L��S{�(o�x�56߅���"
�����Q�� ��r:*����ۃ
����D��	�8�X��Q7l�5�Sl`�A�&�#8��֯�^�-��؊.&b
U�`}:����-��N�X1L8�1��`#���̑NJY5��H�,A�a�R���j!��)0d�i��@1,y���������Q��[3S�veIv{nՊ��d�^"9	-��>�hqL5��M_�/�`<��T��5b8S9N�\Igysjק��2��ޏ�w���@�8��+2%�Y]�^�'�qL$��r�t9���)c ��~��pz!^�M�-��5�i��'a�5ߌʥ�oə���]S0���P`d���;���`��{����w�3�'��u���|��i�3�௕���\�ʕp�����(������<'���EU+�NX|�؀�9�����*(��s���*��G������705����/I?�că���8�P���[�^ѝϖ�?����)��<g�&�g��m���j]p3Q�E@��a"Ym�[��e!��(�x��(���-_P����3N4�<ꨡ��܍��T2����ܟ��SsF�Y�|�����	Hf���*����p-��*||���@�sq���Y~�Ꜷ�gDaU�m ��FC�:�)�`��9b�HDs���n��B[�	��g���*h��VAm�v���]t���&��k����:�v�,Ce)'8����a��~17o_��t�M���F�Ѩ8+{" �K9i*n@��d��W�����q9��#�ۑ6[�[�K��:Ve�(A�	Mk��RO��4��U xi�sbO����&��1��[7����.@2��j�B�� 9<uR1���;.�����Z�'�v�±_g�8u lJ�
��@!�P�M����yG�s������W,BXii'��.�"�X4��d�딢[K�g�
(6nU4mB��x/q3����O�t�{�M��)�xW�xG
����0���x��݈2Wt|�7'�tm�H�Ol�#'�����ҧ�ܺ���(�21'��-��3�pc�E��t�����V��w��0@>  �YeZh�� ��]�I}��ѳ�ߍN�����`{ X ^ZD���~�#t��R�B|&��<�Z��+ix��Pp���ås\?�&'��ܘ~�W���P�#&������v^M����5E�M�\���
Ф���}����eZ�K&���p?�n}F���9�[k�}iB�$F�A���>��i������-ۨW�l��Cޑ ����X�1�Ą�є�Y�M��&!���3F��^TF��ǳ}�;����H��*o:�ʵ��<Oj0 Tb��4o����C(���A�������d7��}n8� Ҵ{�������3aG��(� ո%1Dd\$~�8���~G���l2]z �07�$M�ϝ���� �V���m�O�����hb���A��nYq5�9e d��䓾t��X�O	Z� �#��yښ�sU>�x�j���d3���nq���Y{R��gcn��.��aM���t�0w楻��^�Ƌ��g���Ҷ���E�ŧXby��le��&���B���صi0C�;�|r���<b��R�A��̾�;�L��������!b��R�RgX��\ãOu��S��Jk����2$�?u�0�<F&�g1)��@V5w�������Bݡ�y��;��ҥ��*�^�.�$�r��F�d���E��s��ݮ�[���b͠��C}��ض�vq�b�V��G1%���t%��_���w|'�b�N �ԣ�������Hx����;��\U�	'�L���������l���W��t�����n>�	�)rs�ڽ�I�~���%h�Vf��(-�I2��QM|�v�*��4����3��a����J<y��ԁ��G�G��0�����N�i¹��$���d���5�Pnp��(Z}n%���?�"{B>Gi~����gB(�7��8+��O��Tр�[����圾(����!(���`��¢�V�WR�����}�����k��f��<�v�N{�Ȁ'qh�r
�PZ� i�(�%/-��:l	ݖv�X1�� U� �Z���{�R(�b
��q���4��Ó���`���C%�Ljh�" {�n��C+g��-w<�Fb���e�;`C�[+#.�`�Q���������\P��X�u��=O3���+��a$��S�xQ�9���.�ԁ��Q�z���>�%c�cv���#��5*o&VL:��FqG{7������FHs�xh8,�Ź#o��DdD^8 �A+!vj�eaTl��յq�q(U�D��JS�����Aގ:��jö�t��0�Y�'&)$�P�U�)���X-Ŕ�@��1�G�Q�4gi�O2M���>�:���@�:T�fR}v}����A��&�Q��G>3�!xU�Y���CV�*a��D���1XQ1�k�L�J������?N��s�"E�A�
��/\j�t��L6M��*�q��of��OoZvq\-Ѵ��=!9��g��z$��es1�j���R����=��Z*�Gi#�/|����t`e��,�p�{#[����/�"cbMABM!r
ۅ9�"A$����$�v�鯜|�V�5�)X�g�4��]
��zQ>�N��x��u��a#�.�:&K>#�F*�]�3|hk �-6^<Wi��\�5��W���o�uZ�V�4��{���+��y�κ�#g5��y4D��x<뚽��5��Ҫ�z�VucUl7;���z� �t:ɀҩ�M��#j���=����9��v�gANv�،U<5�I�tJ!n��@�C�[,�9���V|P~�f�	1����6�/Vnv�3�T���3P�%�N�I�BZ h�d��3�
�jO�w[h�U�g�IX՞_:o�e#휷9��L�l(�l��X�1$q��ٲ.5O#�&ш5�B����yr:[>rSQ֒����y���g��N�4R4?�w�������r��=q<�W�\�!�� ;�/biH�~A�;�:�#p���Z��<�C�\B��Εx�*{��ţ��E=^x�WW<&�7f ��4��m¯HV%��'(�A���w���s��������D�ѝUX=}۠������U8�cn �3��.��Qw�)_�Dyq��LG��2Q�����Z�ڪ�,�C��.y����nT��T��u0�������wǤ���/�y��4�Ld��6ԉ�lP�C��p!��K��F����ݾLd��������n$r�hޒ�!� %`�p�pr�� 0�6���83���N����M�J�]��J�ryfE���^xaۚǠfgP�e��3�W�{bѹw�U5&��:�b�� P�$�V��-E,w�}&�gQ�#{;�{\ύ��e���q�Z�2�ZN�;F"1�]�vN����3��\�jD�B�o�ߠ��~r�o�Y\ل'm�מ|�����J'�0[^~X���%�{Jy��t_�y�	պ�c�n 3O��Rn���)��E�0h(�ϩ;)�=�K��m���{'�k���;�2�%�ϊ��X͝=6��?�w*ã�Â^P���bY�f!93{75>rp7�ʘ���
Es�E����m��F�'�s.ݱ鮄���&����74��ɴj���ɩ��� �+��� �y^'�9��B�r�?����йX�Q-���-�x�A�Z
U��!J����%�ğ��gUR(M�i�5�H���g#b!�����f����"�껻���
k�p��,q���3�\b,������P�R��g/�c�t�.wB���:�x��āݥ.����*���&�=eo�v��ϥ!�l�r�zJ�;�1���//u	�'׷ml�9�QrE�x4��B����g%��XM��K�)�P��b���+˔i�Z��]�� ���3	�����h�ޚRj�l�j|k�H�I���=Zq�t�'ǹV�5Hd!�6�,k����72�� �n�%�Oӄ3ԣZҴ�E�eq��G�[Ҹ/Y�D�JQ�M�ɵ/)�5����UȴJ�,ڗ.a $��PN�8�s�c���r�Ė�/e�Y�^U�s�Mǣ4�IR�݉�1�~�L�*�'��c�{#a�/S�v12OvBA��S��t9F���p
��2���^sK��.����<L�S�HP���X�����{�ļ!�P��Kw��9��>a�H^Ū3��ߕ�I���3��Ej��k�JX7�#���]|�_�U3����k�M���ؘA��rNq*�_-�_*~!�9K����p\䀧{.�	�f�����1�&�9�j�3'A�h����V���r�{!��8��v(�-K"�,x��p� <BwP�0zM $�-�Ì��<�d�w�e-��ްe����^f|�k��	0P��ܘ��,��"+���rj��=k��]�k���9KtB���oj˟��j��{�qr:`����&��}��9��'�+���r,�M���/6��l�;��u`Ʉc����In_L�f��}cP���4��ӷ"���tu������+�b��X$>a�2��pf�e(�9W`�LlC 9X�Ɲ���ն_q���$c��z�̭We��"HꇈkV���a�����˅8�O]L=ϣEA<��#�H�?g+��hl�Y�]R�02����_N���hr�(>3%����V�	Z�rN����ƬZGaq�UI�ϩ>`|�Ѣ����i��Vq�+�p��ᜲ�L�����C�i��h(���c��^K��1W�.�N )f��ːd�LG����m|��i �B{������B��؋ÓD������Q�	�$-�gdk7D�,�Gy%'}�w���b�%v/�{xb����;���&�f5���%f���?����;��wg�DѩL���=ٕ����M6q�AYu��(�/)�`*���툜U�=T��dG) ,������kR����(�9u�C���@ݹ��~�q�)�-v��n�|����8� R����뻔��-��d�d�zA���4j�rͼ�&��W����k�⍵��Rv{�$������z�D� �O&F�HB���^�"��L`)Җ��R����T�ؼ6xx<��XP0*�T�/8V\�r�T��� �r��])鵞D��ܰO@c�� ʲ,Zbg�R�u�{L�QW���3|�T��gT�X�6� k��� )U��3J改���(-�SKc�#��a,%���9��g-����i3����[���� ��"��Z�����Y�gX�<
:d�wD���:�_K^�p�����뙤��`@?e�$[��(�����7i�1�dCI����\3��2��O����
s����A�Iӫj�rE��*8?�x�'�rykɖ���%���LHx�-g�(d�%{g[��[�%ʕ�������8�i2���R���C���YJ
R(_��C$��`c��=8$�C9�)��55T��:D���	E�~�1(�e��0$�p	�������M"9_�O�;B��h��
��g� ��,��4�w�ƪR��A�ְ�u�`P��W�I²�9�u���k�*��*�m����!'�����Z~�,�*�Q8��E.��[v�_�*ܷE���j3!����)"9ڭ�k��v)���ِ�<7���ޤO�7��a-�2P
*�ܿ�0Q4��9��lQ��,�piM��@\j���1�E0�.�k_�!c>�	Vf���¨|�-�b�wH����Of5h5����ϴ�<̙չG�S�	{�����"ң�̉8�^��$k��? [���B>���Ȉ����䵨�|�RN�VH,�U ���H#�f'�M�g]���)�jaZ}�h���o@M�y}h���fߙ"��c�Hh��Xk���n��<CY1�6�V��R�Q���ay+!ۣ�,�PL��z��
B���@|��R����=fb�v(U,\�
�����t��į�F���RaKR轩`hdH�T-�"�p����8�S-�W�O�=�)�b���)B����h�i���l��~@�{�˾#� ��sؠ�����$=�u�t��� ��ݰ�ae��,��`�@�}I��N�?��}��ޚ�-��b�=���)����D*�&�d�-�,�����d����&�r3SX3<9qNJSRK[O�V �>�����'��B��P��q���)H� ����	�!?�������9W�gV�ca$�O�D�/a�����H"��xX��L�*1������y��utv7��7fN8Ys��5O����h��ҙ��M- ���?g< G�MV^�V��SC}���$(�oi;��,�a7�\B�o0¦��r����a���9RIg�+Es�i�.�5�) [{�VL?Ȧ��!HuA�_�0"�l$m*���i�r��j�g����hK��qf���⼻m��`����u1_�ލ��CM���
T4�"\��A�T����Y�[/X��T�'m��^١0��]R�µ}��-���d�"Ǖg��Y�Y7mf�<q�S��C1��W�hwiOz'j��-`��N��ʵ�"!p�i0�W�7�����y@��`rf���w���7�T\jQ^Z�oL@�&�'�5����e�&;ܖ�x솛n%,I��*�,I�~:�n�rƏ��]��Z�����$�ӥ�T:p�R�U{����O?��,���j�$9�;o�w�V<�(!A��ؖl�ۀ7�2����-�!w[����r#0��\�ϢS�m7������J���m&��z������!FQh�K��e��=�Q�@��.,���O2;�J�OA��%Q>��8 �Vt��?|ilZ �bwZ�[���������E><F�#��B�j�牽g��=�]�Er��9�HL,<�Wb3ŝ�US�D͹G��ʬ9Є�d~�}�>��J�"���go�6?	G���'�/&�s4����Y� -�� �ԇ
2^�z��9�͎�|?55��E�����x���D��Qe�����2�T�r��(��3��'�'")щ?�e��;廘��̝$��D�����{�n5���PM��h�k�4J��ú�f�$z��R����Ų��w��6ȝG�X �*躵�%!#w�zhC94u��]ߺ��}+U ���&���p�y�F�슂ئ��?����R�s1
����Q��u�5[&l�Dݛ��?����2>�c��5������^�TH�-�|��'~q�J�5g��z��r5�lH(��c�i�ڝ8"��8yڳ��>���4�l�Oq�q�~t��-���<�IΈ5�$�XW��=	���I�
ޖ5s���#&��e�]��$8��(L	��V&AF�/{�߆4>zV�>�+��P�A��_�UE�'	����e��պnA2�*U(���{��?|�V�=#��ѽH�9��@�tT7��.����#�x{4��*UgX��N|A��cty/ah1F��"�LG�2{����uΠ��ڨދ�IM:�;�af���p���ߜ���CV��F���*g�h�-&γtBoC���l�LC^�X�IYL��|S��v��4c� 
f`�q��c�׮����m�a�v�#Ƞ����[�8�����i$�"ǉ͇�#���d��`K�Jj���|��S����� ��w�Jl�S�HZ�-���� ;��d Ad�&���X��H��Dʯ���Y�\�s8ߗ�S'|���) ucqT0�:�Ż�6%]ˣ�?MK�[���WC��z�!�r�C�����Q�ı�&%�N �{�wZ���&������,�e[��7ꗡ�
zcM����MҌ��l�6;P��]WQ�ܨ������D$�z1����<S�O^�#�|3v|�P��a���Pr���g2�e�G�X�r@�~Q�1r��|��q����<��_�W �/��46*�"i1:b �
��"��4�{���?һhp,2��qT��H*��0��&kr s�T6mS����z�1}��?��!ί3�=���H۞�y���[��h�B��Q_bxm���ܰ����>�b�	G朜���#I)��rϵk5�Jwվ���*�����2]aEҕ�e �]p�G�����{�ﳨ[!G�C��";��.��J��V8�l>�n�d4	i#�����\�qvEc�� ��ژ�ߒ�dW�D�)Np�q��Acb�$�Mq2�Ea�����~
��z��f�����?H��h%8��%��=�J������M�\��Yx\B�QGn~Gߧ��i24ް��h���h�	0"*�t���掃���@���O��A]�j��,M9��0M�~2�' ̚�K`&�5�� �:6*�H��������^kP���ac��+:�N�/����������1@g�w�y�dv)�G�rZ��x@F��@��|�Bz��㺸`�� �nLGxh�ǹd��e�jW�����lc]y^`d�&	��p%"}R����F��I`;�1q��pF�l�����5m�p�����%v ���L%&��r�פ��񜻈��>�ď[�;,���:�X5Gd �`4�������P{ �㮬�� ��ܱ��D�1���Wcd/��?�h�ZЀ���bo��r*	��@un0����1��`h�[�{��A8R���@7F�~dH�ɇ���#��us.��͝�Pز��xBW��5��UEϚߞ�iJ��G�V-����{������qV���Z<F�M��ʚ��Ø��s�T�mR����%0\Y�#4���(
ߧ�3�8%�>���hi������r�a����e��P�q�|�W���u�����!R[-?�@XG�N��w~5!��G�bTb�qpx֢:�e����1|��'j���8"��l'��ys��Eȵl�yr��+>1�<Y��A�PO���^�������+���^���z�����g��ꙮ�]��yfCZF"���D)�d���)l�
� p����[�) ���+VC�]L%�I�r�\p'�)��:vIp�5��V�_B-�&�}��bv��/Ry���wC�hZ�u�a�,i�K���eZ����0[�-�`�'�)��F�8���v1T�؋��Ix���)'= :3��Nr]�]Q�,��ܶ���K�'�Q�v�����Guȣz�̾�i�s?�9��^ȏ�Z���ӎ�] �`�BVႇ���{����!��D��R�)��di�U���`�qt8��O��hV����p�Y5��,K���+�����P���?��I�+����zUQ��e^P��j�)Z�3����t���o�&I:x|�����=�� 2��
x������Rs��TE���&��� �m��h<#2*�t�?�>�F1_f�@������j�Єw���:�ju��������X@^e����xF�I�3�J�����X��K�aT@���ַ��'��55	�Cq�$�P��]8�-���W*YރS7$�7<$�＠O���5��06������@�B�G��N��c
צ��O����:� �:�dWR���@�x�br�@� ��;H���M�7q4_�z��`��M$������eɶs�rjXoƚ�vO�զeZ�Q��<��U��u�?Q�p.R��lP�p�R��r5���>o	$���m�oE)�	��[���L;4[c�!-��"��`��5�p୫�T5��U^a��!a"i	�2����8�,�6�1�\c3�����ooE��i��>�GÉ������#�I3Ȏ�{�|���`Z�гg�oz��7h8�4�eq�-0���߿vХ���nW��8Vq��������k��Ě�4���ԗ��pϞ}:���i�<��jh�~2p�	/�����3�+�r�5OJV�Xۚӹ�<�b��P���
��ك����%}��4�l�M^�V�Q,E�]R���y��!^��:�5���;J��� ,��{7zVE��\�4�{v���P����`vS��榤�V��o�0�J��Ӷi/eby(�u� �(�J����S3�ad;�{�����Wv`�����m��Lܣ��/!� ��zj�O��k^%)�P��hg~�׉o*s҆����| � D2ٶ��B�hR�h�7A/T߸,ʷ�6����� ^m�>��#��K� �O_�/GŦ�����F�GǊ��$�JD��TY��95֝d��@�ɞZ��Z5�xQ@g��l��G��Y�q�Ok����$v�_�of����k�q�������P�bg�ڳ�p�^�M�8*!-�
��|�n:<e���W�D�hA�.S���)L��9 {�
�@5栲���	��9���'����`2�Ʒʦ�*j�C,�t�w�T3C��UK��zސ$�9ՔY:w�N�"ӌ�n��k��݇b%�|�/ͣ��-Z�DY�3�	?��J�Qd�)�����~M6
ZA��[�RǨN.[sMnE���mX�<��t6��
����P�}�����0K�5��Z��*���>�U[rCdD��ʉ%���!���DQ:2��?�VcNʣ��x������5Kh���137���T��4�F��@O��@M����B��K����ዄ���jJ�tvV"[}�9��N���Ix���6zՐ������n\~�/�����򷫃����hq�HM[���3@�P��=����v��Bf��!'��r�9Z?�'%?܆`�8X���=�cM2�#��6����Vk-�X��`jA�3(��:��k/^����PI9>z��v�Bv�[��m���q��7��̘!��m��(�/T�����b���io|�����sY,�\yu�D��	`u.��S�J��
�ԫv��;��xUF���� ��7�Iu�
A2Q`�6��eڦ�
�?��/C�8yDy�]}Ǯ�3�³�h��W`1�V���j.�&O�x�F�����$D�����^{�K�G���>=�'r�խ��`J�hzʐ�>1���>/:ʢ���s����
x�b׽��KDsẝ��m^�=�8�Zc5Z߫$��B-B��*�, uC���k���X�V�	Qi�ƅ
��L�~f�~�<}N=�v����i��h"�^^23��h�;�������1��0�v��!E^���$�w�u�?%VU����.��6$m�P)�|
!y�QD���U��߹%#oէ팬�G#��Z�O<wڙ�!�ф+��'b,1�R����	��TU��=S��9��;g&���J7n��ʷZQ4&𢒍�%����댚G��r �Qfٲ`L���  ��������;��,,����6~r�қ�:��xYQ�N��x�'L���F:�'T)*2�*��uBH��c��t��*�s��Əg�u�&��z���m^`��="��t��Ck�A#:�G0�0�����p�,����tf��D�cSՠ|�r�?l�b$�����Έ�K.w��T���|C�ЧY��f�m�H[Wf����	��h�q�~�T��d#'�7f�$�����!�S����+����`K�0��{L���q2�ʻ.c5E�<%<���I`��HTF��[p����#���ᛞ�O�5�ǓՕ��rP��±�k]��D�Dag���S�����/@�R�HɊh0
�Bb��(��k�܋��������oHe[%}��n�#�*)q������@��B����@1q�*�݂)J�*ӄ�H�a�3@?�蔪����W�|j:ş�-�	:d����^z9�!���ҏ���~�3uo/y�b�R&�L �v3��=M�a�˱�+ x�NԊ<��{�"V'�ܧ�B�2kL��o�K���H�a��ጹ�*^��{惜���� Y�����V��/��XXh|͗�I�������)V���g��>0Tje
��܉�\�׏�нT�� ��U��>E(�Ҷ��6*\�1����gR1<20����ARjo&d�n�IU��=B2�'��-��w堏�1)gj�𓦄Ӌ���wK��W��*{w�)E\C��9��%R��-N�y�+w���d��eY$h��!�=���Q�,?]����{.�/6ړ=��*�VՋ`k~ǽDH"m��{\㝽�釿�<����=��X��
��)G�A�9h��R�\D��tn�)�ʍoMc�b{�zo��j�����j���EU�\7��]y--2�Wq��A�����sY˧w����N�����
���ôU��ip9@ �a?�9��I�D�b�����v�)�]Ԋ<�y��8���p�����";�:x)v6�c-���wy�|��;�J<��_]/]���{����ĳ=�>���+�ze;\W�c(/��=��G�'*���d�le$���-ȥ��K����v���,�l�'u[���P�ƅ6�����Y����gj�ϭ������9�^���IB�a�ؕJ�_H����3��;&��W̜Q��3�¿//�延�������R�z�G������V�A,�%/m!{oGZl���W������ /q<�����Yˀ���Ĺ��ux���8����Dc¥�v�YLu'��.,̪ᑴ��(׮�X�\(���ֳ����]��zPf�	�����u+�3ru8:,8�0�m/Ń"�jY�{&n��9�W�ߋ���
�Y�_i�����Mh��1'L^�" ����ª�
�����ӬZj��H LA7��gOd�Ź<�{�6kP�B)�N�Э��� �AKt͈����kw���Q�������-a4r�nu��5-*T�����^�����vJ�[>/�8���9�3ؖ��Т���yD�5=��\n6��+�O�VΈ��U�B@�>��WG�F��1���H�2I�@F�w�i�M�~| �� ���u�b�8�a\*ӎ¢�`w�8��)�\&<�Y�d4w�}o	=�e%�.��l��0h��t��+�wN��܊���45{�O�?EmҚ��B!٭���7�(�A��Íl�qpU���pW�g�P	�dG�j��8.����mF*��`珀�7��
ؙR�|p��c�[0i�*�Ky�x�1�3lb5�~��5�3���P=/4.M���F��ʥAlҎ̟��+��4���M��l/�)ݼϪ�x�� n"��hF��@���V�'�Α	 �̝6����q�V�@��'Q�&s�0f"p�zݘ$���O�X�|~�<4J��n	�+�Τ8�<�p(�Pd[�Q�8��Q�dIu��G��\�K~��"��>�� ����?,��5�z�6KG�V��̕�1c[�t)D���t������+(��O��Z�Ϙ�����u���yG��(G��0.�/c�������cD~��x/�1��s���X�Pb�
���Fo���e���͡���M�����$v�aQ�G��k�h[6K>!��'9�;�I`�i�Bv�/o�b`��!�T����؁M\u{V��H���E?/g��(~�g稒G&xo,���iy��-�X�쳠�tm���~Y=����Hz�eS���l�(n��ጝ��������.���!��7)d�4h7o�W"eq ��G�/��z�Z��$�`ȨE�FsG�gnߨ�,B*�Y^Dg�$(����H�E�Iw�f�VB�ɨ]rLT_� a"�e�l������)���5�yzXD#����Sz��1�G,U2!F�����=��L�fK�y"h�}��B������{��<�|^��.t`I��
�ӳ�����ॺ7=%������ǭR�mœ*b�f<L�[$�T��{|3�z��=��}�YG1s�K��\Y�m^t�3�iu0��Мu��*��{�#ţr�4��jɌ�>cҀ靟-F�/�1��U���������I�Y�e�C�ڟRqe�F�Mjn�����4��$Ы��9H  ����$p1�]�Oѭo;<i>$H�C���S��SN�����yc�	B��}y���,%���y��ӣ�90��]������j��	�R̊��P��W�^��S�W����-8m�Y�����,:lR٘�P���p64��h�p��(U����3��P�i_A<�v� E�� �n�?��GXǕŰ/��ˍSn�m5ީW�$��Q[qGt3���9]d2*ku����p�ý�J���z�����ϯ��6�c��uܵ��`�|̎G&sAct��sh,X�"�RG@����ݻEҭ���B���d.��w$'A���;<��ֵ�Z����c[��dˬjy4ˀ�:!{���܅���/��Ahh�an�
 �a�4�1��~���W�U��_��WLgn�BIYp\.g*}<�.�mB��V�5y6�B�M�	�>�ӕB�	���N8��Xh��)i�]'
��m�&��<���f�*���I�㉀�N���x�����ǥ����ޔ����C��4�p�$�tS��y��1�D�ngִ�%j����^p&���*E({��rC{�!�
�$���iC��x��g���U
�Z� ʷ�v�R?J����V�u��\0����>TR,�/�C����v	M)��~�=�����%��=�|<���/�/h��%�5�p88'��YA�g���r��$���%7�NYo}/�A�y!��Ѥ:�_0����Ȉ?T���������: �n�z��nFC��w<����h���0�+Aո`��|�V���r!�~?[�+��'в��;BXb�n33�hL�^$��>�BzS.�ۇ�"��̵�	<pF���W��d�Us�'���΍��W��hy���vEؗp{��=V�+*]|����I6��X���W�����U]V�\�Xtǰ����93��v����j8��jW���cJ�w|�݅��O�W�ϪjڵL��R��=sON	��;�`�Z<a����ۊ����U�7���w"�����`�W<�í�(,ա�K_c��j|mM 7�:8�TPnϸК��� w��UQ�x�I���O�E��-����	8�巆���<X�ɂt�� �����)�$[�b��q�z^n�)��2�M�c��bw���!P$������*��x��Z�(�Z2�d�O+KJd�G�?4E������û@�f<����"7�N��nb��ЋՐ�"�.fݰa�ƭ���(����h��t닶)���+���w�[��1s��牦2f����������������!� L��!������{����G��-[vL�bM��UE-��r5�@d�o�D �FC�k������ի~�0Os@|T_ΐe�+����+��'�+lu�B�?*���T"U��vh�v=Z^jݭ�g}/���b�<r��zd�HZ�H�K�@*J��VP�l:�{�S$/Jq��(��)�'�����YiC@�v���͙��`I��N}��5ڟ�<y?+&en\L"6�և�4���S���X�M�쬎s�s�Ι#�"G@]��-7�i���9��}����xgY���<E�.�0i�!�n4%o; �a�q���!���e;��	j9��d�T�Œ�-������ëKڏ�Ͳ�js��*�����TF��l�tMm�9}O0�R�߰�&WL�M���y���X�K���D�k�9r#YԔ�?Hry(*#\~_bJ��v�AIѰ��.���Wz"q|�Ղ��#��7���a!��p�O*%C�R���j�}�����oe���h� {��'w��gG�N�AW:��l��N���,�by��i�(�� M���~X� %�g��/��X<�U��hv���,� �K:��t���Y�P=�����ѹ~��P$_n>_!��2��+�"f�O?�-�7��J��m���u�z���������p�%-n5l��	{�Z���e������ܭ��&:>���h:����4�&*�sU�,�qo�` �~��/�UQT��.�^���/!Sb�(��]y\�,�#T���d�Z�`����pR���Qd�G��n	���P�Rr_��P,hA���볆�fi����}#;�#ޞhQR^CD��+�3a�{�	`�Δ����W.M�j^W�������t\QF�I�h���h��%)p�/� �����s�#�1|(�C=QEݲ໹yu��GH?*~���i��ۘ�m�&;�{��q��9tƴ�8W��^��_�*�w5��Chj��`=��o��Zat�7�p���x6KEp���Ϋ��]�êd�'^募����f{C	�c��>�h�
��:�ɾ��4��XVrzè|�~�9A�K�s���?��`:�*u	H���g���2 G5@����ELì�����H����Sp!_t�H��]�%9����=q��P0g�mk���e�p�?,b�ecP7B8�+*`�=i镶�34��μ�;��-����+��vQ�'4�E���f[*�\:�����I��1[Yӗ�W0�c�g#8ur�W�� .©f�j��ݚ`d��^����6��V����������W�5�!�\)�+Y١��,�/�f�؛?D�@_j�A�$kTsЁԈU��T�%���"�;�ױ���~YDֲq�6�����M~�׿����V|S���������Q�����%c�:��7H����Ĵ�T���k�C�}n����Z3�o|u�^Sf����K���\��H_������fS��j)�������DjS��w�6p�IF�#z�sk�!
��C�d�m܅-�>�����<�����D�Ո&��N���ì��v1�+�g5�2���-P�@��ƍc���F���]mʙ�bβ���T�����HPq��n��v��x_��~��Uph�d�F�m��:��c�+dy��
��#:q߳d�o}o�9џ�&H$3)+���Ё�iwTG�A�\Չ)�������m�&�D:FwC��f�������XK��)�lC�Y<ڈ�Ie3�ܜ�~,`>���<��q6�D`U<���_�����z��6�2�#�'�A�=,6#�� Ё`D�t~q>��Ь���FP3�$�R�!�E.3���N������l��	��8)�&ƣ���Z��0+���:��Z���~s�s�oy	�"8!6�_�qny�b��+yƱ���v�]q�d6�� �#j:E�����oCz�nF~ƅ;M������|����b_'�c$�3�	�!yMi@�(^�@�������`�;��V�8�|�������qPՂe@��\��� �̸�^i��
�>�Q�տ w��\�`��ya.��K�`�AL틗p<��;r���`�
,9.��]|��|!k�"��!�YL��ƜX�H���1cؾt�wjw"6vF68���i�`�#�cn��;>�~��A�{��V�%	���s$���G�x8]�`+vԸ0��,� �L�Ru���50�s̏\�t��ɫ[wq��q�D���Ғ"�N1�VڕR��/'t��cNi������6<YԹPX	��w��W��<cҧ��}�6����b��H�:ۥ�h�N>% =�cbP��~_��%Xr�X��^�
{��@�z�Ad��Z]����B��^�H�7�(;i��'$���dQ0V�zT0|8�@�t()�kqpG�hCҼ0�ugЊ��n_[���}���RcB���q&WL2@���y�����N�:��ow���	��G���=����"�eM>�Ô� ��\�}���>���@�����B�H;��@y_Tf�ׇ�`'�����g#��8��x�ҕ����#�+-*�����/�QA0#��b��t����^�W��<nm�L{MGÀ7"`��lM�r�_�����W�4׺��vR%�#�*�y��\��`�[�D�����M��Q	�E�5���/m��7��JU��B�JqN�؍��6��F}��+Y�M��s��=S�}�&��/�j��CGq�����"�{c��ɼ!�W�����$ [=�w>"_\#/}�{4�a3���HAO���B�{�� J>5��cjzbKȄVC����R�Y���o���m��n��h9qp���$kF�]<�c�L�oN���@�j���]��Ek+a`�j�Ho(�����Z ��}����:[U�uZ:ߪ/(�Oe�~޼W� v|�o�R�fu�<pY� 
j�l���
���"m1�+u��+����8k-��4&>|O�GbJ���v5�Ф�&�N�;ej�G�U�]�ֹ�$���6.`()nl՘�ٔaĤ����7�F����,E��Rf�ՎTQ��ʛ�K�Z��l1`p��c��k"�{�a���leO׽�ӝ4����&���?����b����:f6d{m�~(_�w��zt�<��磰���]pM��}����g�;�HCb�k�?�I-�?�G�쒜:�CT̏���9G�5����z�+R� ,�F�݉zd�Y����mh�t�"O�j�a�\ⴡ�O	L�1r��|�[�������:����#�#��z�
�O�~�")��F��P�&J��^3�7��� w�G��g=8d�Z<���r8���˙���<G ����!��JR�{��U"�W�=tS�L�4�N��_�W�C�{�[6L�̾�z�j��r�k=�т����t>[��l^�$��X!܎o�OP�[��������`n�������op,�*pj��G���/;�]̕�B@z�M�{gv��(�A2e��NI�����AոXR�7IV��Md��'����y�5�re{?wt��E�~q��pC���� HTSL�4[�a|�;;&�Z�L��1�U��]��&g����9�Y��;Fo5�< h 2�f�MY��fH��Nu
<�Py�)����,)2H��#�Or���~�O(�d�Cy�՘�{�O���"���>M,&�B�<{��iY�G�"%V��\*���^څ�iI���>��<ً� Pc��(]�o<Eq;b�E����A],�>=e�Ʌ/q���)^�e(w�[��+�8j�D8Í(��y%i�����sF����Nd��
�v�o
W@�$���(�4 �ZA--�w��z]��*�@Fh`QP?L�~�㸱B*�q]?�;�*������i�8�cN#�Ma��X���ro7�����X�o��E�����_�ɿ�Z;6��OO�щD�qE|m���~!JLԧ{��b�[��+%gw����\a�^����X4'�Wa�q�b$	�%��~El],$Ř�1i{+��4y�˄l�HP|;�����7��v��a��I���.�B�X�_��#���b�>��=M��S�;��T8W��s��	�l��u�T�Q�b�j��մ��[�C{DA��;N��N�?��qn|c͹zj����s��rQ�(�?�e� etM��$�#�3�B�0�4EC�C@����ahH�m���F���14��ݬ������1k�j.�Br u��c�e�������.�?6�+���xۅR�P�/�U�|k�ԃ�$(ׅ�qjU+��^��ǯ�p�?�h��r���1ƞ�k/	�#�$H�)���� ?��)�]��j�y[j~���P�U=-.��p�s6Wj��k�1t���ߺ��g�D�@^m������x�qg֑mG���_9�HS$���fve�r\3;	�oe	� kW��)S�lW-x�T�@��m�)���PS�7/��bG��$r�����{�l�74��f)=��^S��OR��2��j�]�q�G\(��еMv��@�\����҈kς	!_����ط}#8l�1vHM���R�ш� ���2���{.���߲�"�oT���#;w�i��(ޢ�a+��.rΔ�&t��&=���ؼ��;_�7�d�cwJ�l�	1�~X��@�6%�`����B���߀Ru���E��e��O>F�=b��N����3x����J��g���>��Ln��o�O�D���Ϳ��*���}/����x�,Hz�x2P\y;��ۗ��ln�!`ׯ$�p�w�{EP<@EJ3���.u��P;�.��cЛ��ٖLH A�L��cB�y��������Q�[��S��4��C�|@�z�??��D0�X[;��gG��%\��n�OSWܺ��bf-��/
-l�`�+�4z�L{2�>��x�m�㝉���^B�?�8�w�����K?9�#~�" �/�!�ϑ�R�_5 �@��<)��Y�o0�\�b�a�Rﭧ���{��C��4�Uq�)xg2
Y<���D>aM#?���S�'��ޯ��BO�B�˕}z��L��;�LC�[@x��*�//�r{H�RC$���&Ǘ�1��d�;f��-o/�u��uQ�[��儿Z�3W��{��6��|��YY�[ܹ���%��ˀ`Cn����9�cG�߇���t��"`��26X(Co?�l��z4��#|C15i��?b�{m�4�����wH�oY��l%<�}Ҕ�0��ԋ8��CC��^��v{�|��<R9�eH�X���n�}U�0}��ɠ�[na���"���l������d 	$���������U���n�H+g* �l!�v�c��0ī�Bs~4�~Q��<Æ@�ş�\(���Ei#E�3YR�m�|o���dٔO��Bh�I
�U�ް�q��j�-b�GW�����v����zX=fV75�V��r��3��tm�ŉ��q���.�Y��F�	��l`Hgh2Hgv�a�א�$�iɆ�B��L���å��1rꬍ\��Q-�m���{y��fۑ�j��`�Rv��K���6���b'��w�� զ����@�>4-����"��S2b|34�!9� �S�33��N��ȞAQ3�t# +���c�,�כ�T#cE��N��a���f0�P�d�po*��P�]\ֽU�5���T��/�-�X��0�R�,�U�U�3�1'N&����_�d�S�s��Dv3���RRqE#�X�[�1���i7v�G��O�Q8{����I#n�$#��K��d�S�f������؃W���"�=��:��wX"͎ �I�.�&�b{����w�Y�>��:��+f��b���Wu��N��3�`���̳}��k�@o^��d��}�Cg!�n�f��B*�Xo)[<��(��,�}v����mn��X���N���ӕ���+�6�0yU�P��+e�oto����~���y��g�h20��OdC�Л�%�G�q%ذ�l)�O�;}IhA�Q�a��8��X������ﴜ}�G�N8��ST�r窷	3���Q��F���3��с �GH��� ��e�M�V� ��ze;�jݬ�F �%6i�n/��Ю�dZ?H�=�e���3�JLly[Թ6�҂u�����@����|R�f)�oS�s��5d�2:l_��J}���-O�����Rq ��A6���R~����	�-b�1A�%�q�eVؖ���C��M���BN	흵���D)B�j%����&΄�XTeo�!Z>�//٫Ў��h&6�:#�0�-�B!�d��3	��Z��=x1�AxU���`+�����T]s��^	���{^5�{���5�wTx~�9/�"J�\� g�9��c@�$G����O���Zse������/_��NqO��̪O!�����:���O�� �M=쮒o��H�b�5<�h�o��H�7�Q7 =�3`9��������ڦXȕ˗��a(���Oh�M�z��Ǖ�i?f�0����"A��\(�#:��5+�w���禶�2�~5o�k�v9?�)L;��앤Fa��dݜ�uKfěMҏL4Ϙ��QC�Pb��q����
��<+7ӷ
�K�^���u���ӻM`�A�������{����c���h;�؎�+��ù.��6Gi[5�ɒe��]���L����j-s�Qy9L�"R��u㱙�ZG�q�0�����O���{����L�Z��wc�tn_�=����vK������5�����ʶۭEV��Hg�l��GXp��0��A��L��6V�k���x���$c�Օu�
��VK�8��o�Ζ#��l)��mP��/����K�K�
2T\����=zDD�6n<��(��W&F$0��Y��a�oT�r,�1���Q#1�����`���2�̫�̪5��$��%l`w�ȱlV��d�1����ߘ�~e�V���-��h�޾��7M��;6Ë��	�<�n��v�ŞTv�J�Pgv���^ţI�������X�y�?$�4�w��;��� ��+��nQ�����|���*�0��>U�Ȼ C���h1���y���--k`�y�� Z��-���}ژs1�O����W1�H?�o�s�P"����@��xȾ�,ę���$A}�I�m[�ҝYA��nER��E�*Xs1W�d�Ҕ��c����rEn�hLK��:З%b�t��P9Y�s@��搉�٦��5�̌4�H�щ4f4p���Qb��y�C�������O�����������;�v�h<�} ��i#���ת!=`�����嶒�w|��A�N�
=�\T�C�2٤����"y��5Q��5
s�U�	�*��h��<�Y��ݱ&����.+O�w�U��=Õ	oh�S׿F]yyfb�o�>W��֯�>t�C��̂���>��9)^A]�Ïb����Q��o�M���k����5b�Z��?݌5K��'=^i���$f�/]�{s�4�l;���+G�a�!������gHr9�|��`T<V���9(r+��ƚB�Z�qK���$����t����f�=�Ji$h?����b����腢�\�&��"���<V3�6 N���eS\�	线s�ˮ���:b ���8i�aVT�}�������ݮ0��'��a`#X�h�z�@�1o��ũ���s����`��A�x�h�Wڔ(����Q�@@�b��b~L��Kp%w��[��lg�H���n�M3ujg�b�9�����G2X8qA��Em�(`��joS�bQ����C.�������&ҳ� 2BtV�h��Te4��΂	���enMޠ��>��l��B;�e"t|�myt����{�*�h�ޏ�_���H�g]��B�oj�¦D���s�����7��]�k���;�bd�D�$�ԄUB�]���G���)�?�\�D�.��HЖj�H���6x�<��1�D���s̛���ǭ�`�r16��̏1�*�6��g;�f^R�d@�b�ms�]�����Y&8p��.���Sj��u�娯'l¿���k�6��� 6;=7Գ��3,ݢ�_�98p�H�0�v2�*��)���L�N/M� �_�Y1��R�.d��.dC6��)�&�� +���8z��ņi}v��Cs'�=��e���!P���ˁ���V���0�(�Ȫf+��wf�U�uAF��NYr�p��i5�Mꐄ:Kc���"j|�U���k ���#��C������ԩ���<�x�Z �%�����C˥���{w-�t+��f~	�:���M����>�In��h��RJ'G���:��?�d�V��SC���`��N\���Ek���� �1�ڑ�4�y�%Y����ແ�ܤ�"J�Q�������(Oݤ�������d6p*c�9���&V�%5�єL�N^�B���.��&$�oo��������^0���F����	�g����>by��i�����q��3L��{��jr�m�|iġ����4N}�����Zʞ�؞���;(~"��g����g��R�9v�ZJ7H�R>�C�Ȇ[�:XW�S6m���@nڭ��j�cfkS��t*֊S�_
�<Yb�zn�n�	��̺���(_���b,n�:�#�|�G��SXX���>� k�҉�qp�3!��GlgTc�_IM}J�^Q�M�6=7_}a�I?����6�s@)pNf�ۮw�w���A?�b����������t���������k�R��3N���n�/gX5��RLd� �Y`�SL��_Lm;��!�#l��Ȭ���>��`�� YSx�=c��N��t_@q5Uv�.I�r>B8��=lt��p���.�܂�u)V]��=1j�1Dͦ�e���Jb`,�X����Xw-gÍ���Fw2`����;X��3��om����Ov&cTU���8*�CZ)���Z�	|z�H���Q(t�O�;���J꟦JA*+�u�Ny�Y9�A�n{L֊{K��דo�����=��K��B��kbJ�e��!0L/|>�T'g�K���[ґ>j~P���/
~��Z�Yr��5��(;����d&��2�L ef��j$vi�ihF�{L��(����4����.��&�5
ez{�;��JO#�e��n�o@�lW�@���_�Q��j�j!���p�`�;�,��>�6WLI��NOeq�N�k��[K�Nh 9s>�R%��� �_���/�ƢZg�w��3j1�Z����x�D�$X���H�'�_}����h���(1�P��-Ӆ��m�/�!��NN҉��	�;�C�U��Uk�0�Y˽W�,��U�(IE|S�+`����(H	^Ұ%FB�4��F�Ƃ�x|õL��p����e,l}��Η�.�A0��䕋�w�5��!�����]#�l-�N7��[f�m^����i�)J��l����)'\�=�szj�)���7k�Q���.C1��)�o�wíD=T�8	�l��m��ףY�oEb����檈�X�ܓ�[����jO1�76��0FU�Զx�tr��C�1��{X�����+��?�p~��`ݯ"�|�B�[?�͉+a��3ZF������X�ݬT�g|�<������_E4Q�M�H������;9�][�x=¶4����2��)pOQJ:CU	��2����w�X�=���}�衞��F �'�}`�;%���S��T��#�f)���&��rr�-�4���l]��!L-��u�&��F��s$^
ǦK�>����_����N�<�2�X��m.R�6��v��v��a��(أL�A��d�!�7+#mȯ��}�X�|}��r���'�Q.�7�A���2��NL�p]��%��U�W��P�T�֧�Щ�#E��c���T��ٳ���ӭ�! ��s��cX�٫����]}����� �"oJ��$���E����  f[u�UDnM������ۨ��,�����\�ގ�]v�4q�y�T����Bo�V�LLw�Q�[lWO���?k��	�&P�%=�iwD�M k�3?r�U��L�g�����M�6,�6 ���}�ų��q�t(A��H�vhY�7bpJd��F+݊�2�� :���8�(iv�T�m�|�xsZ=B��S
˟YZ���N��#���Aq3��~E�}W�rcwX���S�{�x�2��pZ�XT���$�=���j��N&m+,h�36��͠U�(��~���إ�]9	���	)���\�,V���,X*��MVa"�e]Q�5hBCkh�R$�}�V�q�t9PQ��������&I<�+4oN:c:H$�?���a�>�CvZǴ�C~zk��P���sc(e��8.�،��� �2[���ʚ����K��A�C�8�&7�h`p�u*5-n�L�(���;ǥ&��!�]k�^�*{IX�t�w4�`m߷Y�֑�-ǈ�u練K��ۻT�g����+��z��6�gߞ�ۻ��:�Dp���K���p�\�I��Y��(b${B=�IX���E�C���k������1%�X�.��vѧ�#��ij,�]K�������;h��VK_dMR��3q���wǽ&�(6��ã���Ň�=Vj�̊��6v��|LI}�!��Z�g���N����E�����(d�@ ,�q65e�<g]���҅��cl�b���O�,Dш�a�C��<���2��\�� ��ǟ��~٘��Y������Sa����[륪l�͓r>ݔ5EXW.Ra� ��^�>J���e鏬�}}�� ֻO<Q�n�]��(�J�B��m9�zX�f/�Bu���Qh�SG�v\�|�'����ƱU�i��9�a�wI�Gj�zc�ܵ����~�]�w����q�//7�B@� �1$�6����@��WR�t�M_V�����rcV�0�W���4���֪���Y@n��R�t��}�V�q����<^7vԵ�}0�Ũ�(��ؿX��Sɦ���M� ��1-H��*�o}��Ơbpzg����]����qO��=��[�)-�b�Νsи.�hd]�F����S�Km��kc�����W�l�6tVň����l�ċ��PD�6�A+)����*L7��J=-�$�wN�
t ���n�7f���n.�r*��n�D�d��?rD�a�>�!mZ�#�²����&�*2���}1�H�l/��t�
��}|�����F�� ��}���╳���&�t�K�T9y��J��m_(��8���^�{���H {�D3��З������4@������$�Ag�c늂ůg�!�7��v+u�9����3�iV'���2�~5�<M1O��ұ���X$�g��Z#I	�2��!��Q�3@vc��N��ru�ݿ�S�:t�-nK�[(ST���I�x���ͷ�P��~��b͙�ل���d�˃�כF���G_vlv #�0�N������w�
�*��&��B٩���\�-Sj88ZE߳kѕ^ep໭ӣ����ȱ���T9�`#w�ʣ��ni)�;�_M��̰�s���kJ��Y���ۜ�\5&9���xXT�}��=��Q�����߸�(m)����5C��Es��0L����O�����Z���vSz$����Դ��jEC��%<H�?�J�U�~.Nx�(��dH#�9M��ٞ�<z�щ`x�, �HB,�M�u�Ă�M��&q�J�����p����#E�ґ���WwZ�%���"�ԳF����Ձ��_�) v�$�}5�S ��xb��z���'�P�,ɷ����Xu�n�Wڠ�+c!���s�o�+��_za� B�����S+�Å��l �����ޠ.�4�a`%���e����B�w�y��y ��iG������P��='�+���>�(9�}��[�=��Ln�Q�p�N�'\^��d���׋��P��T�M�^/�:��,5��f'��<���Jij��nqq��vk{ф͆�FL�*�㰈ގm�D<�~z��֢��2]����S࠯,�Z8�h1��A~|�u����?��a��W�4w�(�_1�G����u!�B��7��ֲH�R��B7	���.�L57ӆ���Wc��Q���sJc~�!A C��Wd Z2'�e���)(7��������?��/)�f���s0��m#h��e9A��S��x����DN �Ͳ$�Ǵg%��,�������0%�V�K{+�q-������;��H�?�P;A�)�N�P~���p�~t� 6F���S�w�� ��}���Ct���
���X�]��#4����-) �����F�H���[�<���Y�k�r���w/v7���;c]� ~9����<�H��,w��sά�~F�=e�8?9�l�2����C� ���6/��vIАj�u1�\,V�1�h��g�kz�S��NHM(�/����Ƴ��ro��C�����3�L3�!UvudJT]&i���};�
�]���4;��$���8��Trڱ�X�xP|`-*���{	�|L8��2�����tR�����:�n��;����ѵ�]�Uo�B�k��'�_�����g���8و��c��D��yNt:��S� ��,�8��/nhuA��B��O���R㯱>`���M�=Gzc��)�:�dkI���l�J<� ���7܄����N㾺���j3m�j�TlU�oF#�\��@����Ǐ���k��@��#K"Ֆ��� �_��wK�o'4P㟝��h��3�n��9Us	��d��#�)K�}����g���7y~��z����D%�K�=���:��}�89e��]��>�@O���]�@�.7>���FB���mDɻ(`?��ѧE�L[������k��`S;�R�ᓷ�b?A�ϊ�qx�����t�b6�vD^'&{%�T��v�%�Fq&����X��y����w�Gꀟ�#��u�#��J^@]Q��}I�
�$�B�"ֿk��*�A{��\>�E�h%${���J�3�G	�(-��J��6Y2��Љ���z�xZ�
��%�TB��ZR�em�ޤ��;�B�L?�pꔣ'���~� ��T����x��������	���S��<b�l&�C�)�k�L"��QM�r@ � ��A/��s�Y�A�3��&�D��$9����\2ѓWT1��	b�=;آD��3E��V��I���N0�"b|R����MH���no~��!�a��yv���f�炒�'���Hj�*�,<z�a~����9���j$c��&�G��먕�=���m��f�: �x"X�����Z��E��%+�&�Hʡ'@q�(_֟D�^�%U	W�d8*˒��TZ��5��"��YQ���5���pKX���U`ع�/�u� �o����x4H	l��
�Y��#jS��ok˄�78���ŉ�՞���l_>2�ʤ)Ƣ)MW�2Y�c3r��	GE;��RV�p���|Yz҃�g����JnL���3���i�#6�
|i"�Sy��+�p�������G�ʞO��2����??�8�mQ�_���C��^���'ְ-J��86l�f!5�`�1���2�G#�F���}o��5�ϛ�/Z0��h+�-��ﬢ�5��4�]��;�Y�Q�U8�/_�s(�'����_�PyH�F`};Q�8SYGo����Sf���6��@X�I�Bt�T������3��Kza���L�K߯�˘� ����F|�$,��#c9�S�r~��d�s�	[Q4�Vx�$[6�?s�
W]1�T`���o8�����]�	t^������O�uz6� e���M�0��R@� �2iQ Yfd%��h�0�N�t�wo���a	���^����q�V��/�L��t��(���{K�Pud�a�<�5a9r�
 B�}V��-�Q�"W���Zk��0 �-;�������a 8�J�N��P�wҡ�^ړ�#���xљi��lP(h+ZB�O-o ��bA\�Μ�k��F�Et���z����9%��F������jj�A�ay�=�Jb ǲo"r���j��ޚ�kyG$�1q���k��_6/�՞}��H7�+����A��5:}����+�A ��G�]933��A8��C{e痢�2��3UiY5]K�;V�p��޾<Gʊ��n�X���?���,�eQF���Xs )	���1fKѵ�݂<F܂�=6>��M��6Q_�5gߢ@�ww��Й�:ݴ��;�Z5�a�f�nN�k�����)R�j�R��@q�RJ��+R|Z*hb�>��=y3=���?h�2wj����㻅���F�Bn16s0�'�*��ϳO������.M���"r�j�T�%W����M O'�c�T��3��Z$͑p�4*�����v�D`���C �� �{U��>�;��w28��BıdT>{r]Eg���b$eێ���`\�l2Ԙ���`Lu;N�Iw���J������<��D��@/��O�#���)�z��5�CYM�\�f8օ|KK/�q͓/Ŕ�V��?uGqx�2�ud��n���NU�u���E�ѯ��(s��CX��`��H���e��#ݩ�8{�>H��pz��"���W�>,��mvl�!@�����rC�Ɂ�+�So�^�3u��/����A�j'K�Vo1̺��D�A���05���n�1� �7ý��:%��O�� ��*'��H���>8��-�>��2c1��C���_� �0,�ۢV7V���&�ئxsXɹ������1e�E2 �K����ҁ�/hU�-C;�))��b���M�̡�����'�@��@B��0�K(/�~_��'�o�!?W���4��DU�7]y�PFrR�v������Hz`!B��!����<��N9�I���3�W���-�S�] �
�F��z�{�CsL���aL4�[ŲJz�¼�Sp��h��?���c��f��(0D/��ɹ�3�<<��q��$>|�HX�uP���%���Y�P�l*q� �5��[J�uW垑I��5�S6<w}Qf
���||U7����)����¼9�|(��v��VN�dѭ,��;��a(�l����<�(ū���~��H0]��(�e���p�g~OG '(­|�c�:�C�T��t�Yب���?%�%�0z���5��&\RX �(.F��vj�"5���v��<���a��>�kY'�����(���~�䪆J�@W5G��q�%�l$����|��<�g/�	od)�����1,�S~ו�C$W�m���9>Wu+0S���e�?������4�Â�ʶi'��|[�wd|�B�ȓ-x�?���jY.�B����ӼY���&���^W��w��S.�q,"��]�<ސ�ccg3}J�V�9^q��WࠐV���TA�UC&��L�N�t�|7@Oh��[ �Z���#'�1��&����I|Xk���5��p�o�4�d�Qd�wE[p8�tQ����FCAG��V9��%�qJ)<�|����2�6w9���_	�S���m�!M�)�E�s	_/�P9�Il�+z���VK�J�;щs�!c�T��9O����:����"Lkg�iI#���>pQ�"��8����w�߄�|�;3�
d�f��6��4Ov䣌�)�-p~G*Sw'���jTWz"�x=���f��w��χ[�A~�_�@��Q���N��l��d��9q��n0�h��c3�>�TE�7͊����A�!�N������v��z�(����`I��
���5�����-\'�p�iBv.�|���<���zX�x�|RSk:(�|��a�F��^�����,-ۻ�U�Æ���4SYP���l��Y���$�^�Ý�5�t����0#G�(���
�n�~c"�\��o+3'��������p�;�G�߽�?[oX������p�,J�s��P��FjK�u	]��yAz�B�������th��b�7<pΟ����������� �;�����O}`��_�9���;~ҏ8���aw�ԁ[YU�e�X�=�G#�������+��H���}�L;�9��O�M�`��+�k���7~���#�Q�;�:Č]��@/�>恮d��]Jp+kk���7����V�I2��eZ��w�,g��:%�pc�-��x	vw��o��؅0�~f�0`���T��%��/[0|��fJ���7��b�[8o��g�<}�:k���SP�՝��`H�-F���7�4���'��(����dle$�%��;qh�ƨ:b�&�;.1��/��a��O�B=�k,�F�aF�.�}h���u`!UțW�y��KL��U�v�K��1���2�e�������︙:SX��V�f2��l��{O�q��)g��P� � ;
K��0".Y[jS�Wk	�Wa���:.�"q�mo�6v$�8B�pD�i4����1�,<�$�J��:Ǝ���s�� �)"ξ�B�l����gI�H7Ͱ����J�no����Fgr����Fm{���	��w2ih�u*ӳԅ?6E�N}"
=A����Z*K�W𐀘�a�24�y��2o���!J�/(��%ZNZ�6D�[)����Q���$�y�#�D�E�k�+-Ҥ�:ZQ�kcEߪ���6�'��[�I  �odv؎n�#s���U5�~43j�(��JiQc�BW5�=�����1�^�����x���n�E-�'�C���7H�*祜~��ڤc(�ԓ)�C���L��\��lu6�x���K����Ō2�c�xHʳ(ߧ�c�mHG�oݡ\��q��i<� `�
��	:ߤ�FpK��>P����W��<���{?֚�^�6�$x�P�<`����@��>O�	�zzn˔�?0<��i�O#Y�%�2�ܪ��δ�jp#H���x����
AN6�!(��/�S�ި���+}ZE}�0�6��J����x�1���4�bx����I��_%��*�ܖM��������>�yr�d��C��-�.-���	p�D��N��R�G2Rtf{Zs@��S����2�q�+q�O��a�h؇�Q���E\I6#� pGʕ����g���,�c~�&!�r'���.-|�:��ڊ���[�yL���F�5�u�CD�]�N-s.c���S�T`Xe'��Ch�ZR����^lW^�^���|i֕�EB��[��p/϶0�az�C;����𨐔�B�Q��=�<ɰcݷT�Kc�m��on��[R4^O�:��J��(�:�l߄�g���P1���cK���@�	�0�H8MϏ8��}��E��FV�&{l>wU�Q~�>Xj5�����1��˹#f45(���"�~�I/���!��n��et�����Rۈ����i���������I��o�N0Qx��4o��@R"����Ӣ�i�#ế��2C�A��! q�C8͏7	��'�af��M���;$�n�+����ٟ �좘%�oSnd!	�m!��O��/h{}���H#r��X�!`K8�@j��"2�DP�=�-��7x�Y�п�h��Ig����G"��'�j|�����	��f�����RAr��2���eґl翙� �1�0̓̇�9���l@�:c�$���^='�G#���E�k@%P��ɝ��L� �p���ʒ�A��I�j��P�B��:��?p�贆0.���ʥ�Y�},M���8�4^�E���mEb6���sD�� k9�x��������"ZS%�����'dAL�+��A0�v95+�/�8L�-�0���g�!0A޷FR��dus�z�B_�\ϋ�yg�<���O!��Y"_�0�_�zl¿�>�5wM�� ��[�B��f�����r��Jd���j���$�*h���;�8������Z,
�]�	��s{!H�VS=� ��bim�PD��b�'Y�KU���ȏR���K}�{�O&uܠD�b���ó4�+�|�&�7̫̞;-Q�N���`�E h#���0w+mL��H��|���hZ���zM�!c�<���W��N� �,�����t�(q�#�ԥ|G��{	��C��������ưŵ���l�c����i�遐�{�u�l
x�3k���4J���%���:c�d!��m#�Mf|��M�.�+�8/����c�C]�+av�����k�����$"�`p�ҟG�&ϸ9j�[n�,Ĉ�����d,D��$���C�DH�p/�N9�N,���4 ���F� �JY�&�E��6M;���U�]p��á���7������B6���A*�jOP������������"_d�M�?�F)��v�'�KD�{I�`�
�����e:ȱ�1C�!�v<���ğb[	��ܨ�#E�ƣL?�y3���>�tF�Φ�ϋ�F{L\���R&���yBC���#x�&���Y|w\']������vc���Y_���u#ۚ� ����[��&�;�����ah�F��f�t7^CZXb�`�#��^�K��a��2ޭ��㢚	|7��Tx���T�Xn���am�� ��%N§��G|\�y-;v�0�������xz6id��f�V����+6:G��Z/{�ny��jهHK���̍ &�UV�A@���h$�U#W��8p���G��>��U��Š�&��n��
�M:����
�i>���p��ћo3��/����B�7넏��'�7��m8Tf�_�r#?k>g�y�d�CA/`���*x3)���9��P��E"O�غ0 F�jm�B�'�g]�~�@�_�(�Nz]x�ɓ���iٱ����Jd���e�D�"��,h[b��Ħ��O}0�뿽�\JvќQ_�e�����k�EG��6�)1�w*�L1U���E���h�1�8�Y��������Iu�)��D��i	}��L��&�^Acw����ȣ�8,�|�ґJ9��R|'8h��S��<#rq<��m@�����^'��P���i@�0��5�\�| A����11��P�q'6W�v�60�
TB�6���g��Yi�@������đă'��mѡ:9���9L"�[��P�Q.��ݣ�KW&�f!*�����[��gɖ�kk��)j����b59tkW`v�$�<x*���03�<T%�y��"G�Gi�n;v��5�yg/#]@�^�G���=ܬn�mR2+�Z!;p^�{�Gb�CC/�u��2����b�}���I��珖ǹ�T)0/���y,��C���� �����,�#�]lM��t�+$��3HL%g�P�3MlQ����āxq��߯�L���:kX��ji���2��]���UxQ�x�{��5>�ί�tň�
_+��Z�\i�u.�Y�.��՜������3�
+)xQ��\O�%x��"k{e£j�gO���dJQl�������'&�V�vZ�_
��3I_M�s�f�̙���bQy=������؜K�ak}I�,�we�H���-��#Ґy~ѿf��fW��h�~�n%��{���qP@ی�1~�,��u"��J�p	I�k��!��}�8��(���8JH{OR��H�[=l��A3� SҁX,U�j�*8�.��4�e���"�E�3N3�q�"���C���]ϊ�ۡI���jk؄��Jɿ�_�6�Iތ�g=�U�2��ę?�?��]��aq�@
�om� @Q���K˃��z�K|�'X����i���<a�;7`�!+�2�w��s�K��I��f�b�<���#W���)F��I��1gZ���@L#�>.�=���N�S"�1��/,�!E�`�*Y]F��&�!���8#�YY�Mcg���
����3o�'}�S��Ij�h4f�5��}�0�f��{�V���e�j���4��7R�1L:s�WVCF���d�_��d���N	\Ʌ[6���������9K���o�CUf7>a1�o��Wh��?�?+����G�3v
A�=�N�l��^��ݎd�ǔ�L���"OZֻSDB����?�v�����fi~)�סԉs�p*e�3��<Ʌ������	��T�2���k;�O0u1�W�̗�_��ع�4I��	�μ�{�]����y��(�w8����a��-}᪜V���Q�4���z_���.ԅA>J(�w��rҰ�.Ze=�6Ѩ�`v*� � G���L�<���@F�uy�o͞�G�4bw|�AVG�J�=A��J)�*��lͪ<tP/�!NƘ�%����v�Fʱ�,AA��wb���TZ-� ��vЉ��/5'��a����om8�T%|��f)P��hc�'4�.���2D���)���͍$$%ub/�vT�4T�	�w�׆J��^m�N�ߖ9��E�vK�oĕ �z��B=j\�X7\y��wÂf����,06O���3����)8��2OM�T����:+A�5� �l�9ʡSOy�U,����t��f�h�"4�Yٚ#�&�zs���=Oq	0-��³4��x_®D�T������S�o�|q�ĴD���}Y��1�g ���փwϙZ@�HlX%�\������=cJ�-��&�lj���-`���C\M�ߜ�N��m4n���N�m�lK3��KFs*�lZ��+c���Lt���u�R�.���<����f����O��F���g9����Q����qk�T�o��p�_� 'Yhr�b���{28�,���g�{}vfd�:4�Z�KĪ�埭@#�N-|�d�GI�� ��p�	?-a�&r�3L�|I}�B��w"�TI�m@�+��ՊS������:.S��K��P��	������\/��gi�b�t��%�P�>ԡE�>NBER�q)���N��}���u,	Z$R����f(�r���;���v��l�Ȝ��C���@P��]��+�<�MP�,���r7؅X�^?׺��P��_a��MygOu;�?l ��5S덠�8h�AA٦B�;/H &^yJ�{�J �^��D�!�jݺ'{ !���|�w�5sIn���T��kR(�j�vv���5,4�M~�N���$����9#��'��
�����hH���G]D
fMU���U���uap|����������L��2`���=�.V���'��4�TfJL{��2[x;��R�'��CO�DL�j'��i�}��Nq8�/��w���r%%���V��liɞC�hԗ�>w!�@�p2S5X��>���^�?}b���?l�.%�d7b�U�f���ɕ1�F�>�E����,ű鬽i;n���A �ۀ����z!~b�`s��}���&�,l�I�� ��7��C��{�Vy��X��=r�V9\�sm':�68f�u���
�ܱ.��p�ILg���mb{���q?+�`�����#��ƺe@kC���A�Ln�vz�}~TX�&+L��ӸR�;eA�+U���[MW�1Im��N�C�s<�* .�Ԍ]�p��)P8���Z�8��*=�fǭ_����&��qt6��#b��/-�vz�Q�ז+t���*K�s�;��G�����P8IE��w4�J~��k�J�Ё'T��uec)�Mc��j�t��I���eA��ѓ��1!:�r5uf�h�m{<6p��Vlӕ�av�����F����獰Hw��vK0�#Ѿ�����.y�O��V/0��B����k�K��Q���T�h�Q�z���_ ��'���&�AT����_��Ux�;��ǬG&�ݻw���o?�Z�Sv�u�R�د~.�[���Q��< �0-��)�Rp���n��H�����(��	�~�ͬ��!|�}:'�8z�K��Ɣz��ִ�E���=��	;���X��G�O$(蘩J�{ш�R1�fu�\�-}����K�P�6)�{i�]�+z�p��~�y24���;7M��ζ�A���T��N�˻n؈���F��)$�8�����I �FY�����wN����t�v�}���oX�ۍD�L��r�m�\KU���i��Ѳɐm��o�	W��ZO��4�;=�?\�ȇ`1��?�τ۪c͖��%��������D��'q��VR��J�d�4�k��}t�RˈK�@�8깧���p�S��5����ߦ�&Vn�Rؚ����v��9�X�Uҙq�*�DTH0����������ڰ��9�" �Z�R�u2����В�ɹ��M)U���S=j�ͱ �f$�&V�ָ�I�/�H�쥱�
�S'7'�y�cw��^���z��X�K\h�g���x�J��ֿ���Z�K\!����V�~�y��R3����_���_�TQ��<��l\l���p�������C��7�'�H�-
��h3����_�0�K���?�I��k�Ԍ�w��z�ǟ���c�l!W�7)!R�P�Á�ޅv�l���g#+	�Ǧ��! ~K�^>6Y��[ù�����ϙ�Cà���[�}��)��^������u������hzt������l[�[YI�PW���+�޿~��^�_
	��Cqd�[ c�י~�,��d��qD]�|l(�E��%�qV�!���ߝ�bQ%�����D8���$mV�Of�ήI�83���!�8TD������iS��7��u�L	�=p
�:c[�H784��+B�0g��iu�w+<��u��m��52�T���4���B\��v0��nn��
\ ��2/�(�>M�@��;)���SE�{ d�\�tP&��;�3�����u]�6�L͌ߎ��u�k�x�N疙βӺ��� R��Ԣa�QB��>���O�{1:��^1��}�["c� �Y�x�N��b�� #�FcAks?s��qlN�:�_͍Tc����op�\T	�7�&_\��}����RC7'C!� ��ϯ�9IbB���?��f{�Wqث@�nMQ.����V���.C�}j�gV��:E�v2����7Fz!�1��&y��ъf��F\��~�A��1X8��6=�8��@�Y�a2FZ:�R��|��~b�t��q��E��`|OP�%����:���'�+U�f)d�ǝ����y��ƶ�_���pCn4v�9�]��0�*җ��r'�`�`l��>ׄAܳ�<�U��;�4����%	V���`5�I���!dd�}�~{ =I�&���౔���Ez=���B�ۈ�m�Cu��@��h�w����Ex�����;��x<=׎��k5R0���	
	����Ҕ��/�r9+#<6������9��� � ������i�}��&6S�{]5�_S�V� 
��{]���X�W�!���o^Jي��m]��B�c�"�����{�u`�5c7a���l�1���E"<}��|����t�Р��Er��Id�-A�$Yj���D6K��� ����@�ɮmkX�Abz��T��}��,��s#��U��XlT��#���=[�qT���z#��|`�/ �yD�����[@�H� *L�_P�q�����<�M�����9�w�;AҊ+�z�5�`��{�"��`*N8[�V#%��D����7d��CF/A�ŨH�Ғ�m["5���¼����#/��[��C�=겚B���;ʪ�mo����j;��a��ˮ����E���:��ʸ�L��{�$�q�W�U�5�K����C|ru:e��]�x�Eۖ��phm����~�s��- |�ͪm�*�6���!�!z�ɧ�FY&��߱6:(jغQ���C�k�M�� ��'=y��*aTמaa(�݊c��ϛb7V6�b�1�����JĘ��)��pc?4�nq� ����[%l���&�.�G�}|B�}g�o��u�_��
�%3�U�=%gC�k8z����ģ��K��뀞����xN�s"�5���0#������kgV1)M��I9��yJ%���M7�(��HKK+2�+�-fI�pJ ���v˯?z̰��Q�񃄍s�����������O�P�5�}K~FHηu�Z�f�&�H%k��I��\��7�����*����mY�$�{�譤v1�+
H�d{:��g�^���sc� ��ّ����E��F�T�s�<^kR���D-���k���m���A�Rxy`F:n�4/������մһץ�N��z�F`�p5��8���;d�u���\�u/�!�=_�gcpp�GAJx�feqUP�J��8F�L���7=nX��4�P�_{_�R����S���;��2�M�/Ig���4�b9�U�s6g���%�����Xk:=W�Ӹyh�N�Z"�5,Wa1�?0^>{��P��d|�R������Zw�JH�s�ϱ롒��<G��v\�$ō�o���a��jn6�Q)��s(ض���7�~�Xi��������Mlp݇��7�� ��?�t\��n[�}����{��X'L���{��7I�:���1��|o��p܂I_F�<�s����#*@
 �{<)C�\L����Ǹ�=<��Rɗ��"�Ў>@b�o����f-t�c$��@�p��g*�.Hw�^��O@S����q�9b\~��N�z:��{�J�L��&1�������W�u_g�:��Z��#Q����lI�p����*U��#X�����3�""ka��Ψ�s��/Bc�����{��",�p��@�3, W2�����j�f�Z��:"�T�j����;����2���"ñ� �K��3q(w���)@E�I���É���P���8��Qg��'���K����!�d�Oy[.��m�M���*o�#��μٷU?�`�O����x�B�tj�����@�]�7kS�Ać�!p;�8;@@*���8������ބ�,�, �����w�A2�7Fd�bY�ً�o������p���)�>O�Y"qz����A&=�Jyю�\��V��n�I˿���Q����e����Y%}G ^��чf�8� ��UO����B�����5�a�S�hM�<�Ŀ �8�����҂#�i�ӫ�(C�<��k�-_괩x�ngu�E��4�R;L���V-'ϥ��jwZ#�9pY�y=��`r�%������|"G�J6L�"�����bY4f�-��N�>1	�!{���궑m��E�@&���D-sX�bHQ=�PT��e��ubO�o���hb��;��2U���u�i��r�a`�)��<�ڬ�[�xP���+w).+ڑ�N�Q1����r����=Ūf'���ZK�U�W�ٶ�Iŭ��W�ӏ�H�����j���#@J��b{�(9@�1t\�,M�pP�岿�PO������,0$��&��b<��~2N���ɒ�x�@����E�k��y�3i�:�^>��3@V�v�����~�<s��F,&Q�n� v���-�/��*���wF�\�*>/،�:AA�7y���W�}�]�0����ۥ�`�zt���Lc���a��l�ST|�1�x�  �[\���Z��qB�[��~��z�`��2F�V��E���?qJڵq���!���Y�V��|�b��`>�Hp���_�ae��Te(���kX�Ho��e�l���?'�J�ih��v}5e	����˦�,����� ϶�����BZd�'�Z�/gː�c�N~'�xwr�}i�G(P��v,A���r� ���=��E���7�,ȓ)��`5�z�߼ʳ���K	�� 8��}e���w﨏2�h��Dƣ6dP#N��v��}d���$y��`�!s�U��B��zwf_�!1��	�'Ex�w_e��(�z�dG!W3%ǉ�k�BHl��2�聥�ZH�j��kg��j!�z29�&]X:��&��T吏�s�m洮�z�Ǩ��R@ѧ���s�"��	�U؟��n��-��B7�����'2o���B����}}4�����"nҍ,�r(����;��$jL[1۝�ǰ��ٗ'{Ы�]qH��4m4_�A���3b�ސt�/���8�).�Z�-"�|�N2:@����\x�f�Gdw���	�6&��Lݔ��|E_,�]jT��q��e��}Jͮ����k�L�bͳ;�����#�#�����g�v��>�mIA݇���H�>�w�*}��|��x�S��K�nf�UgB~�T�P�I����������!"%�w�.H����HAe~R������:��Q�c�_%J���΀����)ϔl$J��y�"�C�� \��3(½�K|le�(�k�;.��wZ��S�k5����\�<(\9bm`����z�@� �|���c!Jh>����;��f0|	�_c��(�V�˙��s��H�Ssƶ½~�L���:�] ��2;Pdti�6���F��yZ�0ɶڶ?/�:p��F�O�8?̀F�-��l/�+W�8j�Sh�o�RS�ȏ��-����x����.\�8���Α�Y��Eʡݨ0Q$Npw� .4E�lV#�����$3"��~�[���������<�5>��&����(�d_��Ͱ��=�##��g'kp�u�
/��ט���X�6`J�o��e�˫M;|G��y�
DOͶ:����3� ��/�\�.�
3M�?y�2�aM�*�+���4T�\�$ܦ:}KK�~�n��6�.��E� �D=՝M��o�.'���.W�Ƽ���+Z�7���GN�+��?r�l����49��7���þ�����4�ߠ�s��0��Y��ZK@���VKO�� iO��lg�|�4�v�9��#�2�O鏘2�]���2��r�dM�u&��Y-+�����>�2b���șķ���vN����n���q/M��s�,�`�BI�����?\i��pL+zE�`��L4��@#+��G6�^��������1�e'�2�A�cހÐ5>(-���Gi��eW|	n=��(�YU����B��Io.JGH�n5�h�Li���4DnQ�>�@
k�j탎0~Ϸ|�A�k�6��slCࢪ'�1z-�H�K
A�1� &�"a�Q5����:�S2���_E�����j<�gY����(P�v����n�B� ���a]F �%�������[�_JJ� �}u>�_{�h��q�"�|>�@��̺?|��764!������҄�IGأ������ ��!Dm�';��A�/�2k��-�k�����;6��'�Q/� 7<Y��m�E'�<I�Jn<|¤��;����1k�(dP�l���M�!q�_��7�lFNc�u�Ў)4�'��-��JAʪ�r5�D�Z��o ��ƣC���+Ƥ���'���Q^,���"�eIN���۹aN�X����4Ѭ�&�����`Ʊ�0��R� �ř�-��CM�њ��&?����"���tw�� _v� kAN��w�/$���C�2�񀤕Y�פt���Ƕ{`n�`� ��b𷖕���'��?��bp�>h`x,M���b!/t/5�Q��ƬAR\Kw�V"��c���L�h���!�M\�]/��q���g�����7A�6�΅$PV~�g;Z�E5�6\߅z?�LPp���Z����j���Fוo��^nG�JϘ,�h �c(�ۓ���t��4���Wк5�GI1V�,���!�:6�j�ڬه�T�B��)�R`U��?L����&0B�堚�8��Z�!sIk5�E�Ek�:\�X[oK���t���{Uy�)D��#K4{��z�(]�,�!��۝��q�W���Dl\�2Y�d��F��Ո�.��1Szo��A`7�n��b?��QTq��|C'箯R]-�Ld�S����� #�D���t� �؎H���-�n�x��{�}��N�)=�=���]m,v�f����?6�e6��Z @B\�^��w�Y�ޚւF��'�eJ�%h��7�C�-��@.D��s3��{"�;i�b�^���<�̎�E�wmμ�������ϫݞ�J�b��&r?���ѻ73T��t��&�o
�P�a�4a��ϑ×�@�H��8CS��3����?@��pC�!b]�q
��x�kyn�J���H{�������\=�G�Ne��Zƹ��p6"������#|��;NM�
L�'�)4I��K��N�o����޿�
nI��4A�J�=�m�n����4�zrޑc�����i�]����,��~��%��T��W���3��]��JT�WE���rhq��kD4�0�-T��{p2��ݔa��G� P d�R�W��bܧ�AZ4ۗ̅�4c8�͸��S��+ t��<��0�s�V����pi���J���
�Iv�g��?�=���.ξֆ�J��V���	�4*�b��į����WW�ි�G��m�zӄ�_��J�x��u���]JH�U~�����B.���IK��\0�/���!V1�&9�{�ف�{2�.�}y��D{�Ef$L�W�AY��wFҜZv�H���C�"�7w��O��$L�c-��9{�,�r��fw\Iⴟ���t�B� yWV��PcY�����ےW��](�>qٴ�������_�.T�L��xv�x���t���	4Q���ҭ��ʨ8����%h�A����aCܯ 'N���0Z<J���r���g0p�Og6Y��y�{J���~�7�f;Y�l��3�x�\�2b�,������rY���H\!,�;�Y4��
S��T"�-�[9��ދ����K�W��=����U�IWHt����o�9��Yx��?o�Sd��'Q�ᭁI�����q'�x��Q�`���Cԧ@��l�/(tA�v�4g^�ra��h�ʜ�����6_�SD#֟e=�2��;F�w�����3;}��?L�1��=� 4��*�E�W'��I�Pt�l�yᖨe�l���Œ��s�>� �w�J݄_��zd�QK�z�)�ύ֏��&A��9�;�鯭B#Zq�ј�v.s�FR�ȫ���1�b��FTT2�����=��4Cw2�@Y�0���E�.�<E0�C~��8@���������Z=�H���V�T�Wb�$~����\ dGs��J77�������|�p	5y�lP��Zd���g�b���ȧ�y�p���UL�'x������'�$2@�kD�-�@w�:^:B Il�哰Y��/Am�n�&s�tUWP��et��(!NG��Q_d�6��#_����z�m0�s"�˖!�"�ٯ�o�Q´#���;�1	V��r{~�����,�¸!h�8�l��j$�p���3�x���t�:��wB�i+/�����4��8�9%�7Ou��)&�����!C.��
A��v�p@ ʦؖ���O!�S�ݒܒ���jT����W�mA�F]��L���է`5A��K�@��`���@�����jGA%���j�&�� �Z/���|���IW�f��>���
$5�u*ˑ�A�q"�:��ǃ�o|���r/&	����=6�u�:����e��:/Ě����q�V>��P-�������8�q�
y�P�
t�Y��F�9�D�oȵ�_\j�2"���_`�$E�O#�EC�Q?iY����n��~My��,L�m��NF+M^޺���V�*5b��BEP�>ǆ�=K��
�D����4�*$�c�9����_rK���J� �~�B����N'd�!ѯ�����ʧF�4�E�z�WV��~9�Mx�s�g��A�贈;L)�#T>���y
�A�:P�֙��I8օ]��-�k�"��1�E�!`�n>g�=�s���#ccr��l_xX0�^R�)K7bkb+4��1�xwb���`CK2糉�/!������-q�/�B�e����H,�)�Pڸ�0�9B2:M�0�6@U׫�8W�r�9�O��n�������<�҃�������Gv��£'խ&q�vD.�"��9J����N�6���
�gM�s�~� ��n�ژ�º���~��������4VȠ�Ͱ���fz�F�UЂ��5�>���wȕ�G����m�F��ԯ'�k~�%�>���;n�_Q��䘣��<eez����S���7_.D�S�"u,0��d):6L��"���� ��� 3^jy�����޼X��-��h(���)�|?�	Veɻ$�9tl(���|�J��՞�E(�g,���G�
a��@EbA�Ak������p�jZ�Q�y!�e]���$P^-��w��,�)�����>�_����`;o[1#ڧ�Oa�������T�[ke8�I�ϲ�'�Cڈ����O<rr˷�w�Pͫ���.;j��:X��A|�ˉ���I��`�1]_�����0-���ɑBgC	V[�*�# ]'��w.����a�Yt���8Ř��z���5�:+����\L�zE>֐�eדL�_Y��u71&�M0�Y6&��3m#���w_��f��/*gx�����ޅPˣ~�Pלk50��C����:F�����M��&��,�+kv�]�r`����^�$qH	e���[�wҮ��J_����>/հ���G�-hd��:����� �[���b���G��m��g���?�[c<FG��J���h�-�L	�6.��PހD ���)F��LQ�Mr���0�Η��!$=mK�4A�IF��//�?g�1aIWp��ĩ.�+�*hU�+�1F�:).��l\�5�ͺ��������sh[g�h|�Bf
�9��z���F�)G��P%��H8t3��-�����f����[_�Fd1�9~�A�	�a�ax�΍�'�S����0X���X�������?Wa(7t��-���-�/�kK](~��NR3��cKX����Q��Y�`N�pB�Be鋗�Pd�(�~�@ʫ�W���Ê�d�Q�k�������H��0�7��_S?D�-��'IZېE�cJ�;C��������&��X�i>�K�*���҆�45ǯ6ԏ�p��`_'6K�*�O���Izm1���9��Td�%��c���U1)������%)(��H��.d�Cd���z��u��ΰ��۷U]d��D�&�:���XU�D�aU�����i��!�

�},�`c��ش��ܦ}X܏?{zŚL+=
=̇k�Y��$�n���I����]j�a�b�����[SL�O��1Ϙ|(�勴�46��a�BDf5�g}��Hn!Κ��'{�m	�:-�q�eF'��vj�%En��>��c5�����N�(Hh�����ຨW�-��rz��d��f���)r�9w����������F͢��}z|==�ao�- ;
��/իaF�eƈ(���ª��h��D؆9�N�j����y�U3AG�(�	����嘯t�'2w�\5���J��]�����%�Z%�P̬,�+��6�[�`XL����� �+d�%wDa �7�=u���.x|S�nݡ	��v�By�;��a�|*iBX5?��4�.%�8W�E���:�;�Z�6�3�1<c}��k9K���k���t��r��?77'��NH���&��o��x�R|�"�t�x}�{8ڧ[���T;)��u�½i�%�?�0�á$L�Τ��%�Hu2���k�K_ma������A`ڮǿ�͕b�} ��mY��:W�8,Qt'_fb�&�Β��:km��/K������	5:���-ȸ�5B��Zù��f88zg��@�?$�1>c��oH϶��0���r��X7gn�8g�*��8k��S0 /����LR#$��{w���聑p�������%��HY���lpm:�C*r�`�Y�Go�jhlb�"���J�Û^�/�
������fă��>��q{a�9����3�"R���-7�ƟJk@�$�~!,w�Bi�/f�E�fegm��@!E�Ք���-�����h�C�_c�,T��ГiW��F\h�D����hc���Z���_�W@<�R$_c���B��n��.���Di��߂��0�	P�5�b�Y��X�k���;{͡�D";A�U�x����wDTc������ې��"�W��q=U69�5�È_�B��p������ a�V���G��f��Y�8�]{߈RiO�%��n�=����$�p��T.��"t呼LT:!��(�������JءBb`�ړ�YDY��	�7j3�	E�աD�k��3���3.����Uu+�,�ƀ�Vc�SH��6ş���7Cɧ�Js�H+�e��l�1T8��y�8��*(�2�7�Lf�8��L���tsʥc�i��!q�+b��C���(H��1��A^��Ɠ-��i���F�`@mݴ�n~_���z��l�R�nm�\nXM�<��z�-F#h�j`y;~��nш���ibC��/e��x�t����~&'�_x��b���� =��؅E�u��1]sѕ{�C�+��d�:;����ʛ� ��{��N.(����`gJ���yF��[��^	@�*/,2Ė�NԼ)�/[�N���bcKBne�Ak� 2,~t�O�D������q��,�J���e�p*Lf��O�I&�6���$�Ξ�z��׷
���?��#zv�Ҵ4}ZJ�[ =ꃐ �I�.7��f�=G��Y8�ًװ�5?3�������y�{�B��{L�Cs�׿x�����_̛2�Z@�[��\&�:Q�d�y^	�>���,��ԱA�D;-�ʟ�(Ks�\�)�� �u��a��I5ك��I����)M�L�P��g)�K���Lh����;���%Q� N0 ߻�`�..&DrWc�F*���T�Ay��_�o���b��Hfn�ԥȖ۳�6�$�u']D�>�5��oSayNACKJ����ㅀ��{��O�Lx߲�`|з�(��v���W��#�c$p(��W.��L�ҩ�-u~;�ڨ(�.x[$O\9+�d����W��7�fDӴ�Vl wW��+]��K��R���Bu|���e,��y5��E���AH�S���2��&/��"6���\���U
mJ�X� t���jm��"�:PN���\��L���
��OH~��Z>{Bc�}��mA��o�-��oƷ�7X!`�+�.r4,<�Q@��?����$iج�F�&;U����N�1�w O[#��X��\u,��Ѐ�1�(#u��C*�������t��Ue�`_�I>�gK�'����d$�$Ö���,����}!�p���N�_���Z<w�x)1U����^���(���dU�M��'C����P7������8;�|#7
�����
'õ�I%e�$��`C��N�R�K窱!ar11����&˜��2��H�a׃������T���2�-�4Oҧ�Z�Ѝ�i5����SNuz!=W���~
�㳒7�F��/\�kz�m��@���ͩ�
����a����� �y�l��,���%&��Od�2X��Ô��� �:Y!cyɣ3��k��}���x.U�q̪�Y��.I�����1ƺ	S��"۫D
^�7�~�=
(�	�!�J`!LD���nB�=�%�Ayr8�ii.p��	�<�T��Q�@�3'{�)4���^Ƒ�MQ��4O�/����qs��AQ˛�c������D�nYV	��m_}����������X� �w�Z���������iR��ݗv�A�#��wJ���r	�J��9��9�K�w�Ӧ�-�����U�%���ʇ6� �ۻĞ`
B_'�6�tւLe_�u����T����4�$��X�T��O9yC�khlY����B.ߴ���lڎ[���K!�={� �P��s���W�ߠ�*�SӦ+nP�5�Zg.�76��O���6�L�S�L%�d�O�b�D�(���
�d���&���zE*���qh<����N��}�ϳnb�[�Z
p�I�f��'��XG�s�W����$\b+��L�l�j��JO��x��f+���`j�9��� �9�	�2}] ac�Z[բ�z*F����Q4eri,?X�L&�Q�[dC�^��؊�-��Z�NN��Ѭ�4:"�����Ϙa�K��uA� ��#��еK�������+وc��ƛ��	�.cLj���~UE�Fq�Sob�~����uN��c��hP�裿T�(d��2�Yq�R�2>��'�� �p�O��U��]҅A�@k�y7w���>{,����^�=Bޔ�ꍷ"�'����B��ɐ��H�a�z��Z�K�^1�y�8�=�n��>:l8�OP���d(Wa�g�lW�v�p��FU2ͷt�uׯ�ܥ6����}���C��9ݽ�Q� �gB���LU.� K.21�v���"��RRQA~�B��~����!���o����۷�$�ܤ�i+�wSʺV�
�p��`��!�o���H) '�7?v�
�����k�]��i�n�#�����Tó�v�j2ݾmY���. <�q��F��BY� ��~�����^܂u�k6���T�bpǥ�{��ۜ����3+�Ͻ��5�.�Q� NBd�5ك��@�&_��9�O��V��W>�;�_�ۉ�x�G�xm� ����9��P��u~�h@BS}�:Y�z�mk(T�%�]�SC����?�A_�\ �b5����QA�QNb%q�g+<�8��Yǵ\�
2�!B��AaiP*���2����w'�%U��?ݱ�� ��q7tF_�:���0�ZU0u�ځ$���M�ʔ^Z}e
-t?O�E>;�V�e����p�z�MH�M�s�e���D���<#�s�O2��❏�j��o��*��T����M�0���E�4�r��>�&�4���!v�k��xciy�S���+��r�*����b�r�մ�j�zЪ��}tz�v�Gޒ����8��p��4W w~��u�(QP�����$ᆺ�bv�����Щ�b�1:�8s��f� �$<r�F���z����S,����pI�w�"MJg����ϭ}���(��
��h�`���5؏�~)���t������0q�4�8��곚J���V"I�ZۺJ}����V�a����K�6��y�p���O�@�	(V,4����7��y	�}S�4fW�
���>�����Q)�R:��幮��*-z�H��k5!�**��'$Kv���άK�4p;|��ݑ�,?Ɋ5�����Nǿ�d,} ��,E��kw������?'Rmv���B)�!�K�`h�Uˡ��6�|P�� �]/#O�A�6e0��z[)�H��+7PF�q�;Z꾫y7��1�/��j�� 	�7DS|���/L������~ɂ���;��qИc#�����2���A�Y+�*륽Y���,v�pY��.VDud�_8����k�~``bJȪ��Q���J�$��Ԁa�eHY��?�}��!W�1��נ{��3z��� ^b��X���Z��`#�"�����q�T:��#��kp�z���%����՛{_�b�@��FNTh�b�;&m��8֜����Yk�ʑ�����+�㯝4��-?�|���W�ͦ�!��Ҝ�W��x+�	[L9�\���Vَ�<�_`$��]$m��_�a�ph��R��?eH"ܛVn�����v�	����'U�X�����püo%y��j�:�z=�ϳC'v�
ӆ[�y����r{�_`Ӳ�np��*
��G��R� 	}\fvA~%�ve4�r�9M4p@'��1�:���L�n���&�
2lBʤ�Q~�{���"<���G"i�Ɗ��q�-!������Q�u��	�s�n8��A�5~��ܣ�(�!��Gr�».�I�"�6���`>�'����Ϡ�l�hvFu��K`����"�x&Fd쟸8��N#����?��ԥ�ڨ�l�X���&:w�,����&���!?�����r�9~^�%Ѭ��"G�k�"/��`L cV��b�W����#�Q}<�UJ<.tk��]�_G{�#c�_C�ugA��)�]}۳1��5�JRG���t��ɫ��Ie%�3�-�H���Hv�E�[��o��=�:y����8jP���n�/)����&�.��5I#cK	�(Xߡ海�����ꠍz����c�m�}���oE�f�
�c���S:Ĩ�Ly����k�t�Wg]3n#�i*$)�s=?���3�=����nG�q��� ˡJ�Y�S-��_yU G2Ϣ��o��{��u�D(��C��(ov�3BEp��>�`�8�;�t�^��8�K���"���O|��9F�-7R���Q�4|l�|]|G�m�����:9֒���j�Բ8�z�C�*fo����>f�7��m�g�|��� �������=��HH �8zA���ŷ�)4�,�����˒���7td2:��CGL*ǘ��ں��X}sY�{#�Pe�
�6a���M�=!�ms2�Z��^���;��s�i��"�k��&�)Z�`͐V��bp%K�y9g%cE����Nm����'�Ƥ�5r���$a]T�`92�%�2,Z$!Ŭ?P������bHc�PyV<M��s���EX��g)�̏pz�jrr��U_�9O�8,o�>�_5�����a5���E�Ќ���jj؈��w�[Gi��U�a�?A�,��[�S;��s�O��y��Th0LDy6+�n�1�p�d�v^�n�9�/'�W��$��	�'����!m�u�|�a{�����U�9P�K2@�p�\\׃r�����ޗ��͐����n���U2��f	��
(��\4l9l}� �6�tk|�+Ћ+�YC���s���5)m��e�>.���6��_j���J?!O���W��2((�2ɚs>��m~��J�a�/Rog��%�����4 ���o�����F��L$��PWs?��\ɍ�%�������#��xK�U�>�Ņ�v�3�u�'/@�X�i��t:�� �w_؀�V W��6��fմ�>�B����^��u0��g�-�-�}��=/L6Ď�{��~t���0�1���<KCt�C�",��h�a�klxC|�mP�A�^|��t�2_�����ש�GF2Bc�@�ngN�!N��+���68�*��4�/�K�"�O���~��P�%,�_x�VX�^ye<��&����\0�x���ƥ�0e��>����DP.��у�!G$�� ��`f��~S�&y�+"�*�7��Bˊ��!�>it����H�Z8�~�y�;�$`�Б�2?q>�l8S�0E�h��E~=�W�B�֮�Ө����k%���1%tn$,�q��nk�'x�7;뭄҈ćɆQ=��}�pzGq�2��8������u��\ �#�h� X����������N\y�0e�+ȅ�}r��ү��,�"�k���>��7������cz.{F�F�zKI�H��.� �Jr������V����~��
5�Yf��e�7<��L���cV���]�ӏ�4�#X��ԡ&kt��ta��@Iȓ��3D���9�N��\_��-�P�1�ݹO���2=0�	硶0]'�M��.��u���n�٦����R�C0~��1ʤ�WR�<��A�m4ɾ��*���s�D���X/#^4�q��Cjk�P����k��T`g�n���\K\�9��V� nL����7���v�.=>����%8�!-Ӿ���-~*�Pv�oxְB�7��Y'Jgob�e0λ��<W��{���*�Ū��Xq�}ٸ��W��S�#I}��M�go����^$��(�$�>?}�͡M�=��L�{	��ҹ���2�<"�-y$�����68LO�m(��<'��)����%jc1B�'R��e�g(>"��J����ps��T��XmίOᰚ&�Ν��`�3���V�t���U��T��ҹ��Ml�Js^�� �Q�2�wO\�b��L�#��gӆ~�b��!�/ans��>X��|�ۣ�e[���>����i6��6�0c��q��K�	>�m{�*��E��3(~q�ҿ���\q�)2m�#��'��P�Z�=��G6ax��9Ǥ:'���ȽZK���jC�A2�J���8��9�a�tG�"z)E�ڮ�q�~&��%���7_��2�V���}����>�DG��彑�Ս7w��0�y��¯�m4��Y�X\39EJ�����o�y#e����j	���1��}��s6�D@L���	��3c�A?#Yս m��c�&�]�ם)/�V۽�П5���}s6��$�il�VB��$����;������&=E���jG2�C7��p���oN���Z�4���0)4�7��v�,��!�3��H91t�Vſ(ExP��rY��<�Dmz=@q͏�����$=��~E�ilY��j��_�`=���ʭ�̧Y^�%�3ú���<t���(� M�9.�Tl��LVf,������g��7��С�{p1>�^eI�3��W�	����5�i�;��S��l�U0Йly����?���5�	� ��dHd���l��5���ӉM_0�"f�t;@����©P�x�\����������5�̼�:}�#=�(��x��#^�>Z/C�B�x����a����2j�t�2��[*~^�%ϳ�\ٝ�Sr��,B��~��RJ! ~X��M�ߐLk�o����cvU�ͱJ�WA�-�Us�~�3�Ⱦu�97�ǣ�	��	C�v�M��sM��iN�)�:��)����\ց�V�B������Z/�@�{��{��u�5x�ȻKa�����W8�#Ɉ��'�0W_��"A��#�����Ξ��wW�ҽ�.]M�����)���(�N����%�,�r&-��W�T���(�ϳ���<t�7�B����[��,�9��"���B:&"��黸�0�L��E�}\�v����Y��[2ŉ�{X��e��G���[� �d��8��b�'��Cx[��Ħ��q�(|K��u�������c&��k^'��u�ʶ�z��ӿW䢅�G��<���D3U|��۸�[�q�( ��IRSα����Ai�'��?��^�w��1` ����ȗ�C�ܱ�]=��O�~l-<(�ߧ^ZtmiGoӝ���/����k[V������ia�Þ81��U�7ܵ>m��pY�nU��H� m�YVW{�8ڬ�SJq����J�Y@�k�1]�6��|ȁ6��U�α4�$iV��8%��H��x녺X����J�u��|F�t�bpjq~zI䴇���c�������{_1K�������7\-5��0z�`��O��:�U��R�<�������w��
�wF;��9:2�jd
&���&�~����g�I����B���̉���ڝ���碾�qw�"�*�T�A���*c����`�-�kyc������L7�:��|m0��:`t�Yä��{B��2�s����hI�30>盭�c�4���=ۅh���-�R򶮖+)�f[�"���>��)��u�'gXI�p{�~�#A������/����x�u��q���^�)ށ1���j��LU�`3A'�� a����f�H��̃�Wt��n���#N�{Ƈ��,wo_�B�Pn��y@�����ɧ�vѦƕ@�E{O6(v��"X�:e���G�V�l�Z$Ⱥ�-K.Y�|-���P B�-�Y�!D���:�>O����>ј�W���JV�$��1���t3E}����P�ѫt�D�9Y�����-�M���į��_�P�@P�0�����Pc�֍�`/I��T9!�F8C5�¤�F��Dr�I�-O*w�:x������tl_{٦.�d��q墈���'�k��+0�������nx^	^��D�<����E<�H�P�Y�Z�}�KO�֦��R��c���2 t�¸W��ǹ`V��X��ﶾ������ʙ���J��{��}�x����d��xI���1�Ђ��^��uk�a�b��t�%���_2��v��`�m\��-bh��#:�m!$V|3�[�nQO�L@gZJ��� �Rh/e��\g�ŏ�� m����4 '݈�8�ˆ�q�L��;H��\�'�\z�"Fm�8�l�"�4�%����Q@T�H\�+NDtT7ӓn�ti�fqG�)��S+�8����{^�_��&�.���uڲ�`+�Nji�|Y�B�n�=��"e����m��h�K�є�R�6��yn�i,h��2?6�y�yE����(�߀elry��$��V�9�-~����E1�6��K4�u��n��xT}�_���=���2u:PY4#� �wɶ��	M*u�@�	�X���쁩H8���\6b|�Jt���s?�bmN2u��!�S�k��бU���iT�}�+~i�~=@p�+kPџ���<�/���X/h_X\hod,du����zA��&x���V��X����B���#�:���Z�f��e�?�,�lT^����"��di�	����}�k��m��ܿZ $̈���b�#-�4;��ɏ'�:��������.0�>�.$�$�F��z�4!^`=�*s` _T�/�2`��4X3�O���yX�5Al��dmU�Z��_>#f�AU����(��e?$��U�:g.7b�j��Zb5�� ˶<�� {y����ˤ�-��4_����c����QA!�p��T�y����v�.E�ͧ*y]9�-�b����A�	o����ߥ|~���t��,�e<�%UϽ5mN(��&/5b`:�{4�j���)VL�W��!�-���-%��,l｡*���#�hv�&	���9�K-���.}n��(���|}��4��%��*	���L��;� ���31��>���fhb�R�v?�V�:pⒶ!.��?bg䯶W1)�G��
�y��n��i{�>���)Ij���H��S��d�2�VU���h�f��B%��y<���,kǭ8���J�����`W�� Qr�7��|���0d��smL4�<�~l@Cwߜq�WkP���P�] L�a�K�1��f��7Q{�ϱ�����O���Q �N��p^�˾x,���\���tUg�7�j�Y�l������<V����=x1R�a"��%�d`i�� c7
x�֝���ߍ��S�g]��*�����x���SJ�����9�W`��/��Z��,~��,�~�W,�^�T9#���	K�b����^iB��8��g9�m�'0gF���Tw,���v4�6l"������]��X�� ��6���� ׄ�-� �b�K�D����$��`�Sq>Z��i%���������<6�:�(AС�p��C^�"�h@ix�����ӷ\��+�P�]n20�?c�_?5GǛ},�!�ON��D_/͘ߒ�-k#&ǥ�D�I�&6�v��|km)����h*H,��̰=��#^�S��sI%��u�ai/��Y="Ԣ{x�贴2���T�p�cr\.GMf�L�����3�N��yx�8w�n�16��\�,�,ޛ�b�/���K��	`�����*gl ���=h���zQ��&��_7�&�7�k	Ač�0ٻ���.P#���� 1 o=*�F.��Qz��LQ��� ��k��G����i����ʀܥ��.�PaEj���+�|O40l7��+��3��r����O	j�S79���SVU��Ie�(������A�^,�^'~���A�gB+8^L��Pb�F�4ߩаTb�=ȵ��� {���u�Z�����O�ɁX��E{2*������`lC|��,+	�L�e�ش&�߯;MЕz�a�h���B�+oarz拾E���b uy32�޹��Y$V��Yh��D��Nv��)d	E�f��MA�K1������O��,�K�u�W�9c9�s�!�_#�5�.u�&��߉������=gB�M6Ro��c��� ����4u���Nr�O�>������f�c�{ڡ�:N�'*�[M������0~k������8W1
�5����!�����՞���"�Լ r����1��Œ�@����Y��"����qC��EdS��,	>*�f��D6�g|��h0Ta��Q���ߘIoƩ�}�>	%N����U6m�9Ѿ�`�+M��;yt��$/Q�\�,5�4�%E2�0��5,��;�� ��u�8�v~�b��4�L�.��+M�y�s�2*��X�ʦC�(p�m�*��5m������K����M�>j1��:�6��u*p����.��e��/�]����&E,9�?8)�̑\��gH����W���I0#t�|6����_&ȀcČ�|�p�G�ہ^�N$�C���pV��}����5��ƺ�)�3��9fQh�/�z8����pi���Y:��_��]'���E�Dv�<O����{�]ֿݻ՞�sT�m��	�l� �e�o�ai��<{�|���Ó��U1Hu����o🙣z4I �b�1�S�B89,�e��_~D�[��o|WG[�#�fW:�V�G}��"��uR/࿸3a�&:F[w�����E|i	 C5��[�����G<�R�YL�����5��Z鸲�7�iX��4��E�J
�oxz1��C�_.�^������x�P=:7���T��S���E�	_���)�;�H0u�ś��j`s���4���j��F�IVq"fݶ
$s�Q��a,��گ�����u�{j�ar�i�&����^�S~�2���&�7�5�� ��e]��띱�Y�����~�d��g�d�m��/�R8Ӵ���M@�2MZ�j�}����n�.���wɞc�0!U+7˪Ր����X���ȜZ�sN^�E��I�A �T�����@���Hּ�^��9Y����!�`]�˺5���2ʲjG�w?�{1���38���f�i��7��� j���z�b���L&�B2�4,��p���	�s��p���FA��vm�l�}�1lO^�d2n��	"}c�p`Ƨנ��X������f�"Oz2$��f ��y^��KTB�&�~Ǥ�E��5`�����@�ű�Y5�<����z���XZZ���\U�0'��эK�21�.�~�%M*�䋐�Q�3�ļ|�V���sa���=�:�����YuXY-��ݦ��`�=�aj���P��RH%xؕl��C_X�`�Bx��̪ə�o.����Rl ��57}��ՂEY��Wm��*d__�s�X��_6o�?�x��]� Y J<j���x�ߠ_�j�\�<�BP;�cH^R�O4��.��H\��p6�������Ҫ��;�a{�o4�Q�>�-�SP���*C��\6�şV�ՙ�F��A��&}p���H���,`!��a�B��w�:E9�&csJTͼ���Q�W���o��(�V}6e�M����Z>͉?��j;�'YI�Q=�r��_�4裷js�%@Q�֜ӊ�3}K?�}�I�M	K�a��GH�ݸ�Pֽ�ܧϜ�ls��/UB��MC�9�Vx�������>1���ʘL�+�Ӝך�LH�r0���\*R����L4F�<����D�e�ja$w_I��J��;�烬�PT	�S9��$0��]�r�9�l�'�����F��,���j�'���]�X�/�q��a��9����v��068�M�8H��S׋n��1;[�\|7:X�_a=���b+�%t�0LUDR��:*ʘ�%����-�K5�uK� j��?���EYS�£�[-M\�&��o},_�S�2�����Qr���AX�K3�i3I�[����A���ͫ(��
s�7^�f2l��lOTe����qB��٪m���i�>u�Y?�=�� {3Ew�C>�T5�t��l������'j�Ec�χ��,��i{|�+��Oa�K�d/�gᒄ�5;
�f�Do�l[[�BVG��t׭� v�,Zب{c�;5���.k��gel�Y8�9�ʲ#^��^��L��<
�^�+?��Ʃ� ?�c��)|�o󰣊ho�s�/��~e�_>�yf����Qbvy,��9Rr�E3�q�ŝ %Ȋ�p���^�@`�ז)��J}��v����:�r��/��[�P��/���S ��G ^F�fu6	��1��E<�Q���/�$L �Ŀ���uoe-W����9|��PoF'JTt�l2��3[F�δ���(i:7і�y{�|ew���)m�lS��Mb8A�׽��yQ}�^*�Y�R� >��[5��'���#�T:�z��ATz����Ē|,��N��j����>�c/�ǯ����n�1FU�� �*R�s!ҟP
�!�|(G0��҂|��h��o��U�.2O�S	�T�f��5i�.&U{!�ؒ�ܾ���>=���39q�L+.���]�
�0����'��(�z�428�h�Ζ��6�2Ƌ�:?�Yiʣq��^�።F���ܜ�#-V2�o�t��U��Z��!*O���ov>]"z3���e�0��?%a�Ζ �eϬ)$,E}6l������u�a,����
���
hu��W�8!�0d�2�,n���,ﹸme��2�#ߥ��m8�:1r^;�w�����*J��X�G���}z\c���Ș³K"J�β<S����|'��C�Ü�3%�7��<l��ĩK�~],+���	ł��� ��lB]�)��@	��.%t���P��A��[�yB�e9��݄)�D�tJ4A�z�ڳ[�ݳfaJ�V���o\֎����t��0_�'@lؓ�����I��y���F#�ƀ�zu$�pr1�˨�%�gT��d9�	����o0�s�R7+�^	;�<�о��3�6��~�LoR�$&����̝���Q^�,���0E7L'��{�,>��eY���@���`))<h-��	����b���:)�
��g]����M����Bt˶:�fA��Fz�-��X�x�
���%�<m�N��Ěg���h�yO��Ŋ+I�_����^eWiԶ�n��)���F���~�S��f�p܎=�~�+Jc�1-#EZb_U/�a��S��/g�z,��TB젉���IŲ�Tp�G:J�0N�	�-���Y�
�EbޥA��z����K�Q����9�§r۴�Lk�([���E���(N����iJ�����PCjI�si�i��P�/��󝚿!�֓j���q,\��$Y�,�On[b�W��7+�t���+[�%�r`��S�[�m�I����E�č~S�/��PɊ��'y���:KC9�Y�W�z$9^�Q�.EO�UJ�F�}�:��7�Z�\t���|���	"w�vp��|���Lг*���AfM--��S����nƳA8��pA}�_�wF�}�&^�άk*n���L@n�2�b�����C���m���k�� �2��p�nP�/&��ߐMV4g#�ڌ���*��3�(�	��ʸ*��|�|ʟ�- �����x��9�!�g��M
E/н�W ��9�c�� �k�T�x�w�{���W��vS��'�R�(Y̡�Z�/{�[݄E�S4�Q[�X�
����p%��U��I8<�/P� [rI��s�u>]���⭖_^G��vR��ě���vu�� !G �w���H̑8(��� �1��s����@��i��&��Z��f2I}A���_�x���xS���U+�M� �� ����^�*'�|�.��s�ea<D$�s���}�|]���ͱ��	��Ī�D�֜�h�s���#��CZ�
"ټ�Ԁ��(���%�P۔*�&�YB׷�^.dC��!Q�<�7PZٱ_��^�z�/�"u�	}���_I�Mx��������\��S2����m�㐼��I��#�?~����d�b|���x�6s'o@&���{��%RZP_�V���u���h��b�קyG�}+}��.BJW��}		6�-Lb5�7���S�p�Wp�@8c�s`�
GSemu����F!�+_[�à/�t��1<��
O�{Z��������f��	!�$�������f��NM: V�W�B8���$B�x�i��������ERq�EW.�9D.�(?�(C��^���"����\���x��UR����'��V�S�t��9�v��)1�j����I�+L��<�,6�L��xk�c��ƍ�	��Gf�pb{�6I���a����]�:�#yѪQ�n��7.��	�4��]�O�����.�*�P5��d���"�.}GL ��K��˂�? ^�!��S7�P��u�\���Q��Jq��S�'�1�$��]�ϔ>.��­m틼3n�5����S�|Z�ts���ſg;h!mR }g�������sj�ӨA���%����ћEƗg�]o�G^l�ٷ�_��gK gj����~,z���5G���7��~}��s�͇	�p�a�^YR����O����<�S�X�b�)7�r2�f� Z�������sI���)�w�@���Y�Q�X���f�����`-�\�Mg��hG 
`��wO��Ru�;�;�fn_V�շe[,�P{]`/9�e�B�Z���"���۝����[�����x �a[2��=���|sg?�	!xd���"�:Bׯ�B��#�Fa|���y�q8�q����9��AO��+����o��1��� ��ϧW�:�J����a?��MQK�A$�`-�a�EHI�T��n�+ ���fx�QH�Cl|�����-Y�QK�/�]x7�-ҤSQ���[�E�1�"�ݝ P��d8:�AR�� 2���:@ԤC��`�:Q#�8��:�{F�	�x�Ip�LA�|LwgR��H�ȩY\e�e���n��XH�?ZU`��~�j7�����~�&vڢ�IP"��ڱ��8�T�Hl7�v���m�>bd����i������GqZ�1	��+:Yp?*��>����-���K[�O��vޓ��i��:i��b�g���H�����TV����;��D)�%"��UX�e0"��.U@��16���(���X"�¾��@>|
W����w��Yz��s����}��u��Tgvhؿ@b_�����#����T�H��(�u�}ճ���S&��76�IO!j�*n�6o��M�y��9ܒ)�9�0��n>����>ƨ����
L��c�9�x�;Q�\��m5q���W�����B�p�2�D�|�W�m��9���F���\-D�L�l�z^�"(_���u�^*������ph�O��J�(�����٨�1>�-q>z��g�ɐ!t2�����T ܉�JL*P�W�j(b�ڬMZɫN勘v���!�b�=���2��t`�b�Z�\a���Xh�k���?�|���};u_;�{�/ǂ�n��9�5֑�@��� kT�^w)\�:��S6t ����e 1y�3��XBQ[v��� ��:��҂��FE>�O�e�%fK�cIE�躖a!��S쐡Ҿt^qq��!�	����BP��@
�)_O�PC�xK�_>�@h9�9uD��tV���hd�,o�%gaN��9��7�L����Q�n'
bn��?+�A�iH21b�����r�4����� q]m�"e��E�����d����< O��JӉh+�.���J�7�D��X���0S/0$�����Wu}�AU"(�:]*��*��e�>'������;�K᪶�����wB\�yRKh��;%�@;�� :c]�%d�k�E|�&�"@>f�-���͵�+����ڊ��R �����)��jG�~��&��������5%*K{����FT��g�fhB�������8Y�q]|���i�F٘��u ����� ź�����$�uȃ�g�Fo��oolc�_U��Y���E�n�~t��HijRo!�@?Jjh�dl�H-�_�Fgi� '�f;R�F^�[<�L��i%'Y0NF�E� ��Z�R��4�<��[V�����nɰ�q�1.1�gs��뮓����"�3��뱠,L�잢oF�<�U��ߊM0��7:��tj�����T�*,�'=�d�i؂��M}���9�#'��3鲩g���;��d:w����x!�P���2��'���3'W��~�:"-JX��#ۙ�my�nk�Jӳx0��sfh�+F��z��� �U���.J�B�P��$���Yfx�~��������~�1Ϲ;���1%�-E�2v��0lA#���_�_�my�<G����l�.�I��a�E�����g����{���r�V\��{W��Y�%2�n�A�W�=�L�P�򕎺1ŕ@�@D�����\�zL%�WG��
F�le�@�:�д���c�F����Y��X%شh/U������уV�S���/^- ~��G�D���|>y����3���w����4NK9n�3aE�h^�D����i������/8�-�?/��GZ%�ڌ�"MAL���fR�}�OW�1�>�w��'�'��p���@���g�<�S�a8N�8M�F���������g�04�`P3i/�MeV�ڠj&{�k��O��x� �=�Uy-;˹|4�J��.P���	�E��?CMɛ^~���b�Hs�p��To?�x^P+�~��e���a8�v��k�����h�/»��V�[am
�C@��Es/�Nq�P�h�jt/6� l�P+�������A�w�Qk������F���e���Z��\�.a%�;dE1ƶ׉���-dڄ��q�W�&�}�ӷ������*%~hJ��{�K�C+���v��4a`�����C�	��X��k�ZB�֧��ƞI�s�j������L�p�kS=���}#Ȧ�-�P����1���@LSʞ*�̾�.��AEUh I���D�J��gY�o�2:�*��Nf��]��>� ���ȬO��C)�m�;$YG��@��;
7M�ɧz=h���d����#3�X�9<8 )���-t����Ap�!<�v�C9��Ě�w��)��yt0�n=�c0��!��w��9~ټ�g��Kbq��P��rc�ó�J \�
�{��i]�n�����2P�jp�m�Kx��\���m�� +��$BuS3��1,g6������M���J@�+5�މ�c�����G��CI�[�
���vh�����`Ÿ9g�c��^h�OÅnӫy,%kskFs��c�6�FO�	��z}V�)p�����sj Rz��YE1>c[����Ŭs� I�ч�[���%���	����������1�ϵ�L��٪n�	J�V7�0���k(Kڡ�cX�3�9%�;���׀�FTS�`�`�yv�T_�s��H�4Zw��Gm:>PQ�Ϳ�iL�)x�����G�����@�:�����(o��'��E�\���dwNj�<\��}�	H#!�*ݦWԙ"+��j���u��-$��{���
@oD黃�]�P�~��Q=�;������$W�P����y��c�e�v�I1�a9xQ~Ddg��9�]5%�cz+K��[O�Q̭̚W�����O~)�y����vۏ���X^���|ȓ`�5��b�"7�AkO����m?�\��z�9j����pL��kA%\�.Z���	i5�.՚~%g�Jf���n��]���%iD(��R�^Q�7��k���̔��~���D�w;�Q1і��ՌM���	$����幦�2�"-V@T�RǜO��q�SǦ�z���H�=��&�ZX��E����;���r��m�4Z���;�D\���yk�5��}�v��-r�GJPJ)�?�|ES_wLY������#�ո��@�>��Z*�/r�|ￏI�$������|��[J����<q�~K�hѫ��:+>M4E�$����=ͮ0����|z�Yh��e������)����z�B�M'z�c$�����S6�Ǻ�>�(�g��S�9v;sb)�S�����#|��Go�J�!��/��j7f��l����u^�T���ב+�4C�k����hu"���i�e-�H��OU]�r!34���me8���?g��͸]�]��m�6�ᶛ�m�M�%z�Tpt|�!~� ��S��C��M����q-M2ٻ��R��gA����IGϝ7ZLP�ʩre�ԤE�)�
GE"�#�3+5)�2��y�:spR�X�9�!�X]yT�0E3�B��K*�A��n�?�����Z-�6��Nmz� 0��t`�g;-l���kL{vj��:���H��X㇤�K��EC`��`�a���	�C�|E[Q|wKQx����ܴ'���<�z�������&������/6�U�]�/so�(��c��{�s�/𹐈}�5Q�c���"A^��6;jV$ͬ�Q'hqe}q`���ie���zʯ���ؚ�;t@(���V�e΃IU��i^%�s�M�4�1�>m���	�
����*>�oevh#��c�8L��t� @�s�4B�8��vsl_�!�S�8�U����-����!F�'ℽX�;��Ȓpu����F@� ���t&4\T\:��F1V��.�E�kON7�L��&�-x0VH~�p��/�#���Q)%��oCY��l�ɯ����Ժ:�c�]�m<R�+]$��"��T,	�z1��#}S�p&(�=��5�q�^�̀y�b��_��Y��R�.G�)$p�VAT �ߙN�z7c��D����=��>�T���"*@L�����
���]��Tz0�8�;C�wi0�?@6:�7��:cl8Gi����և�*������H���(v$��7������NJ�t�q�H|:��}C��&ݍ/M ��_���	`��� .� ���w&V
!�ﱛ��x(
�
5��)�C�Fۤ;J�	
��{ѻf�#��$&e�R��\
0��;<��$j͕N2邇A� ~^�0�����4v/�ZC�z߻�c�F3��k�������:+_�_D]��<���� [�
�O���[��� Ip��a���OV��y��� z� [þ�M�r΋�{�II�����O�c%S{1%���J�?�|�ym�ܰ�枽>�r*G��r��� I7'ed�����52w4f��x����4щ鼺�JE<�#D&|����!lsĺ]Y!�n�v�EnZG<�$��V��Y�x�PPy��m���ǔ���z,[??����Y#$��ķ}R�]��u����O���>���B&_/H�>�O7.����y���d�����Z���p��Z�7%��gH��g�#Y_J����U�+�pU<&�,��֋����a5x����X�-v�&����ېΐnnIc����De�]��wf٦a�Y}b�8�^��]h�2�r�SBr`�Sz-Tyf�XJ��D��މ����kw���Ap���;i)�����P=|���<���_�c�ta� ?��[�3��6��62�5�N��e�� rQ�1Q�d��o!��/ފ�n�����+��I�4(�u	�q��,6�L���y��LߧJI�o�9�����bk(�z��6<b�L�ˠ���0���U�+YU��""�
p�ct���4E���/0"Y6�0�h�t/�klϧ$)S�~;>i|*�m8��T�OhН�x�T=��,7�-�~=T/w�>�d5g�SF��Nĕg���3�Y2�6�?'T0�=1}ŔKfl�Q"�|�~��\ٛW�Pse�g�R� �~MD��?����s�*�-|YE���<Z�.&Ky;�NI���N����n^��*�qy�|�p�^엀:�?4=�_S��(�N���I\&����"VyJ�+�0�0��y����Z�YL���
���7��p��k9g/^Oz�>D~���[���4�m�.�GZ�U!�b�m!��|G	�
ᔪ��y���Wt)9k5&v-��[_?��v�g��'׵�h�.�[��û�7-�_�TV�1����D!���,������F��HI����{��meÐo%8���-�p��V���B59���WU�]�\�����,���s$�/y6������(\���V�V9{ۙ��&7B���*�r[w4�H
/Z��K@}�!
f\_�fx%' �" �j��V�jq
dNɚ�u����v3Q�֠9����!�9q&��H��W�{W�]�xO�����V��L6�����Ӛ��0P�ҎS �|��mt~lLP�Y
���"ES�v����A�%V��cɰ�zmyO������[��\ϬSI`z����C�ͼ�As��̤����E�֢�X�숆���\�X�{�X��#�o|�G|�� d�x�E�Q��IR�4�V�����62�3ZʢPO���˟LO�X�D2��#�̫��8/w�=�C�T���p����2g�۲�s��~�Mf�[Ex��
3�<�I`Z'!W�_���M��=%=mm�$j��N���R ���0�)�̇��65IǪ�� oVj�YI��!��^�<���ea��S��q90���R��p3*�]I�Q��vW���VK�X�:0Z$��F%g~$,׾�`��D��m[�`s�z�|���MāHG�䎞 8��QS��~o\E��9q�V��I�S�.������(C��m��;t�,a�&SΫ����!��/��aU�`�9��x�0D�Fš�ڞ[���8�e�WR�U,#M�"w jm	 ' ��w�!���.�+�j?��E*Қ��K|-:�|��UO@ˈ[?T���&�!���?������ǢΥ����-�g��N�x���)�_�SP��%�(�siM3����~�$,���<���}ħ��/����̸8����2��p�Ȑ�l��t�9{��Qa+��u��9p͟�jp�٤�lK(��E�˱a�l|�e��N ZY��l:p�+�Ğ�^�tC=��d���hm����u�5�x�v�V�tO�Wr�bn�p��8F5�ڇئ���U1�9�8G��T�$��j1@rɷnw7��|)#�b3�	�����w�2z���у�:�80��ʘ�͐A�;��-s˙�\?v�jW�w�Ew����^���O�;���ز�%cW&&����>�c��3�{�3��=u�&C�g{�5��@�8���յ�)�`��>��m���y�ûc`���'�9�gF����2��@ǆj��.�."�ZYA�,���u���C"�Ǯ+	Ag+6���7A,	,ڝ4������9��d�NqcJ���Ll����k�alhQ���9����X�2�4 u?���T #SQQ�1!��9���d�ҥ�jo�j6F_�P%7p��{�����`�$ٲ�~{T	���
�CD7\�����c�RDql���Y�ռ�%ۨ;�Q'Rp�iѯ'캥�j���"�kz��<-9��"Ʃu!u\��l"�r�rf�:����L����e�y�����OD��Щ �~W_�}ck �H�������i����j�g�����,~�D��#/�4W�؆R@l-�Ԩ Q��'?�X��Î�������ϥF�F�������㒽��!��������F���LM�����qSUX>�Ҟ��m�`��	a
zp�8�N@�L���_��T<7[��d��s}��ڍp~o�.g��'a�AD����x1ׇ\"ŏN�d�u	��-i�OV�3�R����ƃ��ɧb$���A,��N9\�i5ܺs<j<��>C�}�\;�.��d'���5K�a�99ݳ��0�ń�""[5~����H��z�>{B�����lHA���p�Z�MlE������H�J��� �f�|`��T�D
F��#����f�Ё��!�n����cK4����OW�b��ci$3�^�i,�+�e�a�w�$��� ��h�HB��WN��%�䑿�S�,��wݐk�c�h YfF ���ȍc�bk�O[ΥN̵�.	��>����%�4t�׭�n���r)#
8I7~�p�.�d2��H�ť6L<���D-���	;�W@�[���!G�"���A �̹�������+�b���?j��ח���t%ǎ�GGsA�>K���S�7�`�W�k^��S���z�, �+05D����?M~4���e�*�s��vt��V�=���� ����Z8,to.�����շM;n��S=&?�����,YO��>���*�׽��`�����@
�����q�M�@���np�*ش��r6	z�}�M�_γ�Y9��BZd黳�q<;v��ФPYu�O��|�d��n�����Mq��0�lH�ukg��·p@�Me�4~.���%�M�4�#V���I�d�O��z�`�Y��P��1,�,��z�pr,�㔋� ���2���@.�̥��!�G�^��p���?�{���蘾��9�aR�c�h2�tl�)�[�=sU���~�.�N���L��x�L�� '�w�f��^m����Jܧ`��Jo"�������_�S�H�gӰ�~�&p��7S������٭��cl~�M���Z��!�A���n�G�.�
�M���GPٔ �D��Y%������(tpq�����?�,F\� �gK��d�7�u��ס�����?��}�K�$������o	2�d�u,���dm�i�����5�Ω�S1p��Q�e�9Ĳ�n����wp=�T��4qb�Ix������o��,_�^h��x��Iy5EE�{���ų�� )Ys�M��i`�~+�y60�Z��ۀ'p�L	R�cU�o�BT�om���c9��Ys�E�������P�u-(A�_�[$E���mZ�"Ȧ1��
���D.����l�\��RT�$	x�d�v�� 3�2���S��aJ�}�tT�ﲘ�)��.vH�KPO���~D��TjW"U��oi���4Q�����<0�'�.w+-;<ף��(?%����>�A��B��A����W�M(�<q�/-	�i8M��@��!�M�iO�[��J0�p�/M̯���֮.���>�+W�O�rzτ�,�ʎ�PX���Q�P�|qfY�(���ߑR�u��[s����n)�,ޕ]ہ��1�h|-��'T!"@��"m+�}�s�ٴ��n�3Ӷ>�v�e}�];�����L����2`[X7X{�c�����Ub�~����P��tn�m�C������BA=qB�����0)�V�ipmץ-��W}�P���L�)~��������[V�&�[IRߋ��.��������:���4_�;����b-��ܙ �����}1�o�;��� P��Bw�s/u��A��3�wk�{(G���8�Os��)�ϙ�s���d٩��S4G�ĸM�E�co��J��W����(+����m.O$߁'0΢6�ڮI�����)��|w�~a��7M�Kdu�1��%y���,i�J���
����%�����-�⎿s���uZ��]�����s��|ܲ�����L~T���! qU"~Z��� �m�����ٌ���&�KY����������se�@�b4�id��wA�t�},m/	�r�ի�م������}Q������dr�PlA
aZ���*���1�<ۗ��lϓN &JC�yt}��6����E<{��-$��(Z��:GĒ�pB�f��d~�T_@���\���J��eC�Cw>��/�U�B�=���B��[����W"�`���:1]��ˊ|��pHU�����W�D��\��	��=�?���ɨ���q�N��,Z-����+P�B�!��z{di�2Wu�XKE ��#Y.'Q�©�c)�p��-�(޺|����שR1�g��a�|�SȃO	ᜂXvd|.���a�r��5ȧ6�?LT��-y�J�t9�ʚ_.N�����)*>O�9
�
�4��i��+��6:�90����h�b\ZK<� /�AO�S�\�{��C��cK����<ª�1��0]�4Z�;�V��G�*��Jr_]��23�H@U���1>[ �w���=\X΢y|��0AV�P���(i��qc�*s�Y��$5Ҹsl�6�be�0���5:�����\��J���U׌����
M5B#�Ax��|���P�X�M1j�{�d�jA����	m��ο�]����81�A{�E�)dJ3�A0�?���<GuW�0!��Ρ��� �3�c�}�p��B`��Sw�&:�F*��������Д���tN���Q54h��C�D8�^�ա��y���֙�f9�
y'<�K�P��9�M�̬/=MB�C��࿍��G��DO79�����R�����H[D(�)��Ы�*�.x��H�tH̤\���,���D14�G���B��2f��+�ϓ�{�4C�`�y5��zֱk/f��GO�UL��d�7�K�)�mV��|.�	��k/�����E��O��J��#M�.+j�)����g��h:��A#�N�LWY�peu������^�ٴ�]0s���Ae~�-G��x`��=9"M�&��)I��aʢ�!^Do����o$i�Ez��`2�����I��.L:j(��{�c�	���u��y
��e.nt���+z|*��F@3��?>K#�e�]�QF���r�"���v̾{}�38��qp�}m)�w �G��B������\�4�_�CZէ��X��  ��m�6�7���^�|��F�Q!�De���
�g�G��Pi��	�b�<ꂇ�^�pۨ@�9c^*��j:>��N�	[@�����K�N�b&��}�v�J�5ڕ4
���v�H���FyH�L�3� �ȕV�A�+|y����ܲ�+����.�������v^�7�� Ѥ�v9t��; %M+��thE�] ��J���WO�30��/^�Ώ �~߸+/�S��a���3�/�}<��iI�w��g@IVZ��	���t�D�IF|m�j�!%�0���:���y?G��Wr��<�/!^�Y�MמO_-�5!��L��:�>�x���d�u��ؖ_'O1�{�O��J�kӉi=r�M��! J2�"��2�sX���'�.>/Pp9+E}�^��<BfN����W�����A��p
��%���|�F�ILB�Lo�MQ.����~rE�V3?q��:1�{*�����>�� w@_@�����֒�/n��f�h�<)�{!`��P�� ��52�)uн����H��7px7H9�������a1��-Aɴ��%��	;Ip������.<L?��>���Ǣ �U�F�&��J|EE�9�
.G�#f��ݠ�ca�!j���C_/6%���D�R��y�_;� C8�_xj�Zl_9�>�����g�rʣpb�z+��!����Z\�s;=����j钬"n�Rpٮp���:��p\I�4ud��	���Ӳ���(y�})Ru�?y!�n��>4R�k��z��K��O=���B��E�C\��`R����1�<�)����ɍ���"%�S�}RO�u��VSl�8m����^�#~��.�\���UT�+Q�)��auH.�R�|?�7�ҊYvf/.�)��d�Ov	��L(/�Cl݇o3���Km-�y����Q��g
���V����-���U�k��y��ܠy�)�a���蘠R��ʚ$���Wfxd�S�.ݚh��ĳw�665׾yQ�t��{���j���58���ӏ!l�gm����ђ����_�7xg�������a����(��{�8�"�m1Q>���0�7�&��K�ѡOw�Q������Mg�0Ա��lrf�Q_��������S����ȔW�K����b��J÷��t�[X�В#�K�Mr�`��ʬV���`	��K�(��/.����'bQzG���Gv8Z qKm�zg��ps�*Ccqʋ���O��N���U��MtF���&���r=G��Uk�Ubn��q8���V�+��*|��]4��(*.N����5ݾG�$�'��4���':.w
(�j�̈O���Gf#�U]&M�]��9-t�Y��wjӷdӛI�Wi�Dh_)�@��B���|��"���FP`�� ��#L���/�'g;�I5��F��M���P�7��L��Ճ9��%G ��:f��3w���vB���g� oCcj�������)ʠб�>��̴��L�6��U��┤+:��y�tKX>:/҄�͜�^M�u���L�i5�T�p��j���l*��j�]��Dݼ;�d��@���w]*3m3Gr���[�0�����b����m^������g£ Y��*T�J���e�2S�Uz��[�Qk���*��^f��ۥtN�0)U�y�Dl���B?�^�|!��]W����t�F1#0{�z�)C���(>�;B���&�3S�����m�AGV�5����D���@�'�>�q�vtHZ���
��8r�i��j��N ;��e�����p,W~N�b����s[6k1p0�8�t�db�d7��In<�O�,��N�g����>���������$b�N�!^տ��T���.���]4i�ζ��#���E���c�<���16��荚:H%����� �� �����{�q
G�g}]>I35NX���T��ƚ�Ű�t�M�om��W�����|�����v.���Ρ��G���Ș�������Q_�M`�fF`Lۿ����ω��+Iپ4�cWF��
��RII����S7�9�
��`���6%��w��N�R]!��
�)�UEqI`܃~�]uh�e2���GX���ȁ.}kU�-�sКP�V�f��R�.�������c�=��7; 3b�5p-��j�ݤ������&ОY��K�wNVz��C������a{e�b0Ռ&�ǵ��a��tgf����[N`RyE�Q��E&�r#1Ɲ����x��lZs��-GT�a������(nT���D5���F9Ђ&�@�w����<w�W��9wo��+X�o��$L���f���52Ё�.F6(����7��Ek�Zq�$�� {���ȉ"0V��f d�uԍ��@0s�7�򄧧��pz'd��`���U�o�x�WՊv�|�|Ϊ��B�O-���������5[��ۺ�^L$��I+TҔFDJŻ-|�H��^�z��˪y�_t\� ����@�x�ּ�3���CY�``?�vM}�����5w�Bøp��Q e��u�v���/�̿ʓ�ū�BXO��l+C��s��|��Ǟ��B��� ^��(k
�m"����̓v�/<�P��	��H�e��)e�\eu��C���-�5��f�^^g���h
�~<�%�-�}�f�[g�{1R����>��}D�-m���h����ǠF������Cu��'����W��t�<��B��Av�U,�f4F(�vP�,����R��Mtl��w\�yi���� �os�C�_���k�����	��b�3�f�E��21�vp�B{�b�ˀf3�5<�C��;P���7�2u�61���{�8�k`J��dK�$�u$tc���<G,���f�$o�iE=1�gm�J�ASAo��1���")�Br�����`����E���Bm���Xx(yB��Tl6D,
� � �?6h�o�<{�(���fi/��* =xp�����m �#�Qr�(�\aԜk,JaA�~����O���i��]uOL�E�SV��B���j&'�G�()���:�d��Pd�d��r�r�6��� �G��ۅ��c}��+�L�Q���=`��cG�e���Nn:������$F�b�0:�*����$�>�!6ӗ�TlKT
�����쫼��=����cH�U��ɾ,"IV�ܟi��Ad˰Gk��8��o~�)�QI�/�`E���3ʠ��+J���t�t]����?/w<�R��D�	 �9�D=jo�]�dq
�܈$�����d x.��L)����%�h�^�c	cAڡ�'p�tIވ*gܖKw]��s�3H�Y[�)8v�F>��m��B5�-tAt�G���S w=aކ.Bk"{p�L�w��=^��8��W���Q���e���pFN
���@Mz�[��'����ݳN�ݻ涷c�j��k|=�����Q�����S�E����z1�YtD�O�O��5�nY��w�S��+�}fB��o����c�#)4	�|� ��l��넏�֯K-�כ�`���Y�t�,� �8��r�E�X�Ǉ��Zf�k�LcN+�"d$i�KU�[�WL�ǜ�ѵ�]��#<k	rN�Y��<�y��H� ���d�Ԏ��+��L�4�R�%ya�oz+x���J(ݳ��O-��@v�J�ˑ�O���T#FI��i�X�\L:���&�p\T����?po�>�T���T�|� ��P��r{���z�3��
v���)b�Z6�ѕz��ySE��L9�}$08�8����(�o�|NWi	w�)B�d�ǢC�D�8r�}Q�(���-�v�u������痹"�t���YF�)�%�?mז5��1�$
�i�ymU4E�#��?���Q���R�O�ȿ ��BG�1�qZ�(��<���Spma���U�$c_:��o�DMl��ښ�[=�#
�H9Vas���0����>���(�R1��ꀓq�%�1�<�;����W)���!S�nR�$}B���0F�/��84�+r��@Oe�t�i@��B?�.f�U��#1��)��cY9O&~�j�ÁX�Q��A⻿�)vl|:*�ǘ�u��1 s�z@�{�h⫩K#�K��%�I�&[g��P��בy}?�w�_�M9�t��0P�!���\�p�l���x�Hq�65Im���i��0��L���R�J`Ws�^�'�R�.�?�h(Anr$u��Ӌ�A�vB"�e�K���T��!W
:yQ��LȎ�y�0��1�j���o�佥i*�W�|��S����}\�P�d��XI���#��E�ň'M�J�Vo�1��9�B$�t�$
���ZM��ƽ{�qo����j�O��-���']ط��`�,�'$��;-1/*��Wk+�B�7����mF���fl1�x�w%�@�y�J�'+��������G5q�n؏$ ��Cڼ'�B}��(��K3hШl��,�!E
�c��L9|g	μ���$�!��ڴr����IJ�9��i�b��0"bUo\��c�@�5Kw�I�6��d��(�~����ȧ�\��$��'ȅ/��xW�����wE*5<퓪��a�_$/E���M�D����&���)(mX�,�AߋgU��o��xKg|�}��t�A��!��c�\l@c����t£�%�!�pǳ�Z_2���j"D�B��ͪ?:w�n��?^fL�ʑ5�h,~.2_�8�`N{���K��C`X'"� �T��D�5�w���gj	O�CZ���s��3�˙�p5v�>�Z-����G�#?��X���x�qa�]�]W�<5�Cc�͐M:%R��fc�0 Xy`���������l��e3ȳ�b�T(�!j��������=~��[�Y�����y���G���&�(�g�^k�A�Ѿ��NӰ� �7s���(m9b&��E"ٷ�m�^�wao��&��p���$� �p�T?k�Qf��F[�z6�ݏL�&�;#;�<zQ.���!����M�;�?sJĒ �<��|;w,�(�ii���7)y�eHɔǦ-�1�"��$h��������+��v�I{��A~�`Q����5ZP�wff;Uѕ�x�U���v�p��t�r��Z�p��+�nO��������qVd;�ɪ���%B��<�#y4��LU�;K{J~v�"���u���J�c
�N+RF��O �Q":�M�E�ϯ�=ك�hG�� ��S:'��g/B-B߶�WDVh�������S��ظ6,Y��U�,�%pd�)��C��l�?��ïȔ�˂
ն�B�^;����B
w�
䣦�藑&� Hu��/l^��=:f��:e�����J9R��f?��ڡ��#ٳ$����XC���ܸ��(>��\�E�e��[pd��(|
��v���P���Al�,.Zk��~��b01�ݡXZ�\�7��O^ysNU ���H�~m��1�zp�5�w�d �QZ��n��y*�O��ȁ�o�U�T"�ؖÄ��`��3j�n�S�<��,Lڕ�%����m��	>�a!L�ܳ��ͩj�ܙ�v�����c2�3� ��6O;����&5�'�hΒ��\#�f�)��gMň����O3���Q�O��� �q�\�b�� �n���*�	�
v�dsA�n���{��H�|�~��	�b�۲���M��AFK��m:�&�dp@�w.�.��}�p���',=�@,y���u�ץ��e�c|ĳ��Y=�K��8�#;ܑ�3LW7}��I\戻�,w�%��H�.�t�E�=D����:Ҵ���bc��$ s��A"]��3�'<��FCޅ�e�F达�.7ƫ ^��樹����,PS��8�Ж`��Z;��@�.[���ްf�:���ux��0��p��oX��!�G?� `,�1N�e��=f�}P������5V͵�R.������8�v�"��Bu[�E��E7���v �.Aa�7:�V�玆��S}����&����|iŧCy����lzZ3�ES7���ñ������5�l��{G\�t��x�eٽ�-�A�F��&��D}���'d�|�� �s�ӓ�,���,�u)Y1+ݨ��w�ևI�rr��s;�]U>�^]$�Ǝ��v�>�~�ȎF�^L_�F�l-�ԁ@��c'��O4B���T	����\@[��Ga��]������I�b=��`g<���&��f�D7SO|B���W�d��6���˥��=�$ ����w�˷��l�7�tʯ�J7�r�@��9�K�h��ܣ�:J���i`�*s�>g��k
%����9�������7�������O�ǿ9�O5�i�y�����/�e��P�W�9vm�i�Ia@��j=���%���(BDL��#����,��'�11Q�Ù��#���w	_�����"�{��8�[�ee������1�J�y
�^�s����jw?����g6�|��ϪPwb,�	�~�ev��_��$6Na^�Q$^�0�Mi���ȩ ���2D
����
D@٭�V�D<�\�^R��P�XV�q���!iFk�p���\{��y�.)!X�W
�"�V"�5�uYp�ѫr��DJ�\St���7�ᄿ~!�N��+��j߄
;D��i��6R��Y�`��ky��K�RI�sx�W!�����4��|x�0a��F�&�������p�ù�*fOLSxW��[�D&z��݇�۲k�I��9�;��s7,�Ҩ�,K`*�ߥApw��hq���sw�  ���Q&uҠ���T��!6v�5{��&wh�PlҊD�X�Y��a�g�N��Gi��:��U"c�8����T�c�LV`LӸL�L	��p���`\��3ņ0A*�2� z�[k���0�ݱ 9T�HM�����@n��\�}��N������U՟�'�,�c�_BpK���z��o����V_��"U��
A<�PV���������C�T�Ϧ��o�F6���:�kv76�>�R�ci༤��'Z��I�?��d��.�0<��	����4�ՕAU����%���6)�i:Ԍ�~�6�������3���"���=��DB��-���Ҷ�:��u���hA�!	ͤ#[mE0(x���z�|��Ǭz���e}u�I3#P,d�n,看���x�?yM�����B���Ut���}��C�c�t(;�C����U?�n�P��i��M��K%��W���Г,�����R�5i_�3�۪����Tɺ����&.2~?�z�|f1��
$[�9L���$�o�mUwK�=�+ݼa��T3�����*���c))��n��P�tK���[�B�ߏ�^V�ǹ�oHY���ڶ"�?���ՔvfT��ck0叺ߞ$�>f�-��Z��Fa�5E*��]��Iڸ��	����2����e+�ܓ���Ǻ���<}�P={T�=L��a���v�;v�9/�wkI+_����ə��?`��Ze9-R������1!8m��4}LbP�>A��T=��))q:��HDB�K,T���.:��@�����5��5!�o�z�\?t�y�S���б�ةA�?g�5�g����Lt��ݟ�VZJ4�K���P�H���bM�$�C��ԅͱ����j�Tޚ�}][�]�ZZ< �m�v���e�k1�܀�{��l����p�����>4��'V�}�9�u�:)-��u t���Q�d"Fl�/���;�^�N�Å�<����L/��z�;��\}֓�y�;L|��T+���N굍%�U��Bs�ej�J@�x��d���	;��(@����|�Js%0�D�P��s)�9y����
�w�M�����s���U���.DZ�r�˕�Y���T���Sy�]��yF�F|mܟ���:6�b`ϺLI�\\���~������Rg8h�Eɤ�2���K*_S`#ru5D{u���撃��!&UJ[��` ���B�D�V߱��`�#��E�������Cr�n�9ˑ���~��䇩}���y�7��lm�RW��%Ro����c�v���i�:���xJA1Я�d䘕��.����5�q�8� V�;��]��	j/Y�N4]��;|�ZW����Ӹq���qﱉM₫ƽ�y�x؟k����Ưr��b���{�!�.�h�����d"��u���k8T�V�:&��'�!�9ʧl��d�#8t�H��y���*��L�	Z/�9�zn$��p}g~�rgQ�c��.�:BW3���i����@�$2Vb�+	]%�*� 6%��t]M��Mn2C��(=iu�5��`G��Z�>:�<�L?!���>�x�uX�CUZ�o�V��]�wu�t��,g�܁����>����)F����<�2��4��??�
9�8(N�יɵ�\��	��S}��\ 	&�y'��m\��O|_gy<c,���`�ޏ�^�}X��0����%*��Cő��'A�Nҥ:�=rG�vl�Ox�d��0��@���'��}�Y�E��&�4Z�A=	:� '�$�+w�*�B�.�Oُ�H�!5h�;���j�f����~�Jp� ��"Bv(�i�hW IkP�����
	�_UW�no�`�RK�Dזl|/�t�y=I����ٍA�*�:�|� [�	��3hȣ[�5���Y"��M�6��Q=2:'��q�7�"vޗ������"��{���O*u�>C�}����!R�����e���17�y���]6>m��k���%���T�7�;(�M�F$�@G5�_�;J����z�u�7��E�x>��T\����r�{�}rl�~ԕ-C۠���r	����wͧ�`�����1"���M�4��1Q�9��{�e$3u�������d!��S��`��#�B-���I�l�9�,	���٦�|���1\J߻yaC#�a�a+�r�:ܾG;���G�o݊�Y�(���p�s��R��N���M�:���������IE�Ɯyu�\C���B�7�z��%�Ԧ�~�IdWO |H��zS+���&{��+�|��v��]Nx0b�ҭ*kߢ�䳙2J!)��<��A8�%q�Р�؀݂��'nKU�1��X
0�E9�Es[��i�j�t�t�Oh3;�_Z���ى1�3�_�[l��/��a���e�Munɵ1B/��.�̭�S�������_1�//l�2��?��ƫ���SRF��$6D�"ٳl���+�_A<z�Y�Tę[�yǘ*����Ѱ���܉Co[���Go���0.�m�A �f�\/]���������{�6�<Ő�u�+;Tlɜޣ^��R�r���HN�}1Ti�c7�D��':m3d[@;ƂH�e��,�D�&k{�9O���jh%fI�]�_4 �K��5�Q�*�3V���lQQ�4 ��L��>��P���<4ps�)�(j�qx��U3�ni+-�+��4���n#C��*��	JF�m
�	:Q�另�{�
�ߦ�(��2���B��wO�%�i���hهb0*�����u��m`��8
�^�=�+2@'q�׏7���UZ��u�c����A�o@#����������?|�W��n�9��"C#��y�s�WLIޅ)X�=HC�i%S��`�B@6yگ�z>��OʯDkh�%���C�vRTE�6`��	��2"����OAU.��V����X�ƈ��ꙧEt��$�\�o�z��2�x��u���%�W�0V/��@��Qw>�Z,�0��f
�_ �L�ػ0|uy�����B/@��%�ʟ�iA�r~�KH�����%Q�������k��c��!��^Oip�>��ՓEҺ��v]��Q��4��ڟ�n]qla̎!�" �=��8�J�d� 3�q����ׁ����:$?*!��O2���l*��&L�j|u_��N}ܸ_<@٢`�0�A<��>�SK���a��	O�r�Q��K5��  �tZ�P�?^X����� <a�pH< ��m2<��p�1�F���r��t��i�-%q]ƲՔNb��HM,�"�V��{�dz��4e���\���Z����Z]z��޻�J��� �J.��-�u"�#�*�V�ǋ��l���gY����!\#3a1� ��Y\��H2���|Uo)��"��� }�?L�;�q<�o�_���C�I��z��a]~��-��#y:D�3	�&�_x�No�2�{��$��Ҍcf��m IX0~��;�,;{h}�C�@k"�~����l�@I�J�%��z~��Me���v��h�њ��j�-
��\�/��w�6�8_������;mOي�I���HY��d���W�l��<P;J��$������1�8��E����[����}H&U����Wz��`<'�D7{�A���FZ(�9�x�c=���b]��l�Z�]�\
>�"�7���m&�Gu�C_�?��!����X'1'�t��-lP4M陀��7~/��o#ht�!�I�$��=�����$�iO��oNg��<�l(ȥ��fW�.�U���~7e����Xb��e�T�_�7E�8/�12��\�4Xۤ��޳�s�F�ɝ�B�ښ7O������1&�Q+!�xe����no�!�zf6�D���j/���R ]g���끺�-�wFQp�&�~'Q>��#���:���
�%$��������#�2�L���1HR{������Y(+�&�rңR`\V9��[����O{Jg��P�v w{�b�
��[Mr�9ۀ	���u�ǚ�]����X=��A߼.�aEs�sm�4>*�kđ�3���/��u���ԗ|6�D8:��E�l�Ђj��D���*s����+۫�1�q����r��RE��T�+��H��UB�8�$�������'�5]]:�D�	���[H\ݔѓI���ϷF4Q�� �[�y�L"��|!�g�&7��r� �����3�[��\�(�0
�� ���I<�t�U��m�<�NB��opjw�@�\�V�>c_��([��D3]�I�F	���>��X�56�eWX�V.�y�?�L�:�G�����2�m�w�6q	X�JSI�Ҕ6�hΠ�A"�,��[����MI����R�#:ԏz�?��߽��Cj~�7��b���u�=�,¤���4aq��������n��I �AO���P�g���Np�4��~��`�f�1�Լ�-e5�� wg&])�8�W���O�p/5(����a�N��9�5��R����������EC�Zt@�J��!���X0�_���2��+�*g8�Pp�o��{Sdj���9R�]��*��6���bfbtN�:Mb���-
���k�T�hk�ш��:k+�1ֵV4� x Ձ�O	c��M���M��8�	�'��HVP_Kz��ι䯝��r��U���]feu��i\��O����E��n	��?�����S7@�)JI"�%@z|��H�,j��a������r�Qecpa�BҶ�i�Rӭ|����zp{���Z }�1ي����KM��jxY|�P�R�(�RJҞuz�ͤ;9�{�B��@l^����^��.� �£%lXq,&����;Tc�{,CYOs��H��A{s�s�Gh�,b�7���Q���7�
�O����[�v�!���4E/��Z��ՠE�_��6Q8>��.���8F�;�7�,[@:�F^J� ��v��D�Г3��T�8d���tJA������S�v:x�<�Ɍ�7�B�(+! �W�p]j?}����@^�n��]cR� ߈ ����*Ā��g(ʿ ��d0�}�]�5�p�QƯ���>�o�z�����t�*��l��az�CV����%'�Z�� ��7��o}�i�.���M_�� 3)�����s���'X��~��n@A�%C���7D��C*=�y|	�
�$l�B*4��s<x$1PȄR�RAx��c�ⅉ�iA�%�nl����ů�*��B��9�D�6�L<��}�a��'��YVo[��(��E��+]����3�m�W���"�%�֚�]�
���Þ8�=+F���c��R<o�=�o�˱��n��Z% .W�e�TRo���)�Q��� �U�4�i~��N[�EZji$����Ϛ���@a���߀�+������z^?L�I�/HT5�5�������֪�+�	3y��V,R�����U��p�ty���a�Rv|�"U��G7.y���*��'S���4a��y�K�n��b�=�D+�9d��k �H2���Y�0��n��#@��U��2a,����h����`�x����j��B�=~�H�#��G?LQb���"j4�0���; �c��&����&���L�xs/��u���x��mkϩ�c]ʔL����ø�չ`���P2�^7����[L ����j߽ԭ<���e��`�@Y4�3k�k(b�_��I��;h��'��?���'K��At����eC��a��`}���9��/��X���rnZ��P~�`�>�k8�k)x�b|eOd�î��'U��E���	� �@�\;���?����*�]g�{��y�����Bj�V��&V��!sn����a݂��u���o�פ�?�2Z��A��s�=FͤH�R߰!����)���Y�jЕ	#<�8q���$���V�eK�R���M��%f##O�B�����Z�Fh������3.����ؽF�3�S|�� �>	E�:0�� {0����e���R|����`c���I?�ԅjҋ�#�������L�߳U�q�����o&6)Ҭ��; �pC|LO�7v%	��>j���<�X:�0��t��EC���-�hX8~���jb���֛f�t1��5b
��D�<� ͕d	I��.)��4�>��w�=�l�~?h���dm�,c�~���u:��Z��?#\w"���_%%��pG�@���L6��=�ݕ^؄.�֍!`vㄭ~���K��Ђ+e�������mݼ«e�+�ɶ�d�ŭ��<A����a��H��z�%	,e����Sh�Ǖ�����P���a�l����E�/ФN��7�N�ʓ���,��T>�6h� 鍲���E��'���=�`o҇z��nK����jCDa\��>�h��DԀ����©�������TVVt�#wݏ����9�S���˛��s�n�=Y�zEF_4oȻGs�6*-���Td��F]{�������5�9`^ԛG�-�E�[P"�B�5���$B�:����_]�'%�)��O��Jz��������0Rp����?4�f�ڀ�h2cATSy��u�)U$�E��ǚ����]�W%�Ѹ��(�nD�-�Gæ�%c�#˒��w䔹&.K 2m��&���B�����Qʿwn�)`�І<|�.P��]�8��H�߇�%R`7e5�ľl��
�v ��\��1�#��r�'�t�﨣n"r���F��>�ۅ�sg�I�¡M���y�L���ח���OqS��:���Rz\�����ċ��k�F}.�J�O��$A������æ��]�.��*GQ�]ICkx��aa���̧C�T@���J �NZd�P��Vn ��z{��igaS�J����0O�E�qo�q�	熭v@OG5�rpa��-���^�J�� �%?�&�*:�{z�N	��"R��|ؼٚ�u�V(�JO�m/����s����%b����/t�����U%'{��c2���U8[�l�b���[�_ݰ?��-�3M(~��n�8���7^=70��M�e���	5��QL�*KP%�aA���ry4d��/� ���{ �����m��\j�ߥ˧U�q�8�:�	R��.x�����G���2
E��N�]��z���	)���}�m����bu��/�6�{gX�����xf��_v��)䒄?M��SE�8*�h��p�����ʙ�a�>�������-�*�}��>w#�=s�ɫZ�S��dy���B[��	JP�W�s����9<"/����kTW%Om��\�R2��e���%��t��+S�[~b �;���QM�Y��lm�2pW��U�ul56|dI�./IQ`�E��\������ո�����Y�L_��MGJr!+D�C�t�E��3|1~AM��lN4�ކ��ap�h2|-pb��'�G3��=��M?96S���*Q gg>Ύ���.��\�:��J��~"$�X�d5�t���ւ'��s�K�6���:Z+�,�X��[��Y�;0+=�\u�uHE��s�z����lH;a=Şx��0���R!Q��g���/n2C���SS�z������~����?���@D�����]�}V<!���t����Y�Q�)��
xX/Ljq_� �q�2��:_~,�����-�z���r�������M����E�E���rN`%�%[9�ʌ�2t�ԑ���R�2WUc.}W�u.���/\��(���%P���_w���O�>��hQ��7c��?����*���-��c���q�p���$�|��]���04��'�O��j�����mW���-6pXA.Y�?�B	����m�w�j�F`�z���ИHD���1���{W�]���"J�6o����
�&���H�e@���R���y��g��LV����U�8��C�@)� B*ŗ�M� Pau.6����5'�xN7U���c�h��Ƣ8;�X��Xe�a��#��s��������q��3�4����j� 7��0G=D�I���+J4���p���H��L;��0�������)n9"�jYB��k��񑷂}j��&^�ka�O��>�$A֨_ a�je�<��e_{�-!P��WF��r����(0�6L!���ĥ�`�$�`*��!ϊF6ǲch�zU4��N&#�}>�i��x�>��n]d��H>�}}�hΩ�<W���\/ě�99����r}9�%��ɛ}Z�-BlgA�f{��z^�t�M_���=�ա�0�M*���lk"oXc��t�_�}ȡ�?�7���3���<�=�
���f��
�	�=χ��ս`k��!��R6�9��U#B��/-�ȡ�]��j��,�#,7��$*.���b�5�Ss���Z����^C�lA��c���Vk��{�{=�;> W��-'�@�<�P�xϨ�
m�P_yc���	k�V��s�@r8B����s��n��`3�l����o6�+
��X��T��z}��?v���;?|C�K`fבc����%����1�ɿ��p�t�0�D�)�RS�佴/���F1��W>X�B/�{��O�_�O�7���,�^�2O��η���o��4�J�����{�b����J�	��4�8��H��B�>t�xd����WXѿ(�$0<dz6hث�@?�p]�	_6�!UxS�7�5+��{ o���қ��]9�Ġ+0�oTo̘��ݓ�(�Q�1��;M�ݽd�7u̯�:_���Ȍ�J=~�n&�-�H&r�O���2�h*�a�rbi|`���<d��Dt�,���P��V��Ud��Z�_��0w鄬���p;��;�C��΃@t��9ƣ�!3']T�W�uW6:y�j�����{�P2�5VԢ��,��~��ꢹ�_ 5���@$$���6$��]Nh>)��=K�X��"�4�6˰L��{���>���#M0� m|�iۊ2�FM֝_�m�õ:�cP�z�h^�8,vv˫�TѠ���3 ����z�bM�w�������/`��x�]����B��{�������^OS�~�������'M��*G���!�qp��LZwN���l#���y�D�`���xclPY�kǴ�� �T���ϣ �һ����%��$"S�RAUq��`W�ڔiW����&�%@��Y+�&�}�TƠ�����/e�<Jέxi�m\Ab@H��1j&e���&T�Ss��(��W��wK(Q5��W�mUM
�
ze7{��8�~�d3�{;�/k�T�G�m5�O����������[׀��jRg���q͋ QK������豄I��CEO�Y�_��g�"���m�-�L!~!J'lk���k�x;��׈���X�=�K㜟�
ߖ�2
���S��9a`�g�r	"���X�k4t�ݑx��1&??��Xbsư�nN�n�"��|G����Γ��p�$�Tڤ��x{t��M͆��G�R��f�B��Ç�-��Y�錮���K�4����t�1g?�2���nK�u(���a�㤰�;>�)���}�b��8p1;��	_���}���t��
�O�D�U4�	�(u������|��oһ��ٙ$*堧
����T!�`�ꎯ�&0.&������.�'-�40A�3�βT�\G
��V������yP=��؏=(ojb#s�"U�K���3����y�";�/<���l^2{�5� J2�_�I��0�#�����.�O��}�G��FS�%J�;,���8k�1�R���.6S��?�?��N����"�І�m���h϶���GnF>m�DBo��Y1�ם�^��	��[)���j>u�O�m�{<2B��}#�c�Uz�j����?�qE<�D�&�F�~�$Y]�,�Tk�l�1v3�[�?��~�P@�+����>�L���9��V���Ċ��4�S�)-�b��%�{񉺷ԗ��kCz���,�ܘ�[��5����JoT,����N�Z�t"�?�&��f83�u~a\p5���x68W�`���q��Y7��[�Sg���>z�Nk@����Ŧ�b%G�"/��~[���t�s�YƗ]`|6����y`7��j�2��A���i��p1�1k.kUv�5�fwD��G��R�J5lg�h�ځ9�<��~ԩ�-�ߨ�p�%o�i3XʀΈa�����YUVIgsIC�s 漓��Ŏ��vJ
Л�*,C�p��ƨ��;G��Wh��,K�V����1A���M �IAY�	��ز]����G�L �4Ms ^Z=_3�"�-@!��:�Ȝ��bP��R&� �G+����p/���\��{��]��3� �h�6�gN@A��I.�:���JN����g<cҊ��۔)c�:��HGݦ��<}sc�c���) ���4Že� -{{GZ|ޓk�OL�1�YQ���UZ/�;N�n����ۨ?b�5-���R=�����ëB�Ĩ	p� [�R<���6��D��]�9���H�� ��D]����讨� VոU>����Ai$��*�J��Q� �2��m�:��^<1J��M��af���m6�4�y��0�Rv�\�{fG>5]jK4BC<!�x
�1��m!���Ydd����r,��ϊ�������r��T�.�s*]162��x,� d�q�^z�Xʎ1p�;;S��*�MO?�ҿrf��bM���ID����r��柩��*ǂ�Y3�V�U�IeL�ʡo)�0Aq�{��m�m��ܹ�I]��=�<f�
Hۘ�����O�B�i���P���.��&KdKX��:�	o�����Y�|��Z�(�o�O็|����?\�? Y��*BP�U��a.zM9LHs�9�SH��Z�	p*�1�m>�x��:��r�.տ�Q}�;�\Ճռ�0h�@�Kѽ0|���OO�3|GT7}H���3��	�i$�S��=r ���7�ЍDGƠE�G��h�uU����1�}'��y�[����k��}�j����$��n���>��	$޴�)0R�a�����J����~V�t�|mZ\:^rR���jAB��%���ߐT��9�Vh0��Y/��	t'����L�u���^��G'��v�ᴝ>Ab�3's)#���$~`9%����Bm
��թmU:U ��3|�����"�i}�L�*XkIi��n����l��{�^�b��O�6,Y\Z�M�[X4��BR�TU���v��~�7����
�F\F�l�����r �[�up�V�b�vB�����(O��!��D&>�n�-��PTY?�-\R�-�7��5�#���L��;L%�Ц�mdOB
�1�i�k��떴�9�Fy��1�t�U)���a�В^§�OZצ'"{��3���XEG���"������W+���r����x�U�J���R:�[Qqw\"�C�.��؝ȁ4��o���&q���+���7c�+ a��Q�6仩��ܹ�8���`K�������9)�ͭi\K�n+�����a��H��|]��Q�B��:S_���y|а��ż�<?O	nΐ��7��d�-���R�p�q9�Pe
z(J���Go�Ҍ�
N����kL����=XG��.W�~�����sG����U���M+?�^	��x��N�2]�x���Ut��y3(���<C��Xo#-�HIQ~
M�.>[����� �2S6��6ʤ��Wf�/�һ�ߠkJ�gͽ�?�rTՉ�䙎MN>س����`41��J��x�t<e~f&���E�{����;�3����*A���)�%�H�� aآ"Z��'X�9݋�H�0O�v`�E�I�X�|j�_0�Zkz�?gU���|g������:L:(%p@���q�R�J�ykQ�c4N~+�XS<39R�����>��d���{�����
V�0.�L���tl�mc�R@����c
��-�g��o�-��aY��G�y!���r� �]5����a\�ܔYH�'>�b��$Ih�xy;��; �FҾ�o^�I�h%�ݚ��M4=��A�
>�@���PU7�_e|SwP�v��:�N���yw!�S���X��l9ā��m�H�=���5��*�\�:�4nLڎr��'�����-2L�`�+<2_-�?�~���>f������xGq�aD�P-��z�N}~�)3��H.���sR\�S�*X��Gˠ��A�&���l�Ѝ�;Q�{#yW�2�U6j,d��M~c�N) ��S__�94�[af����|����si	i�{k(4;�0��߃0�\eb���YK��VM�/K��'t�*¢e͏��� ·F��|d���*�Eן�-*1�b����f<����a�oߞ�y{�|;�$��ס����y(W��?V���MC����=C�̤9wAWN9I�N����*2Ϛ uq��PX7���/NǴa��֔���M�}9%��D��ٺd��Љ�Byq�M�63��R5�	+��3ؚI��a1)�k�.��8�W/�7Nib����C�8�Ľ��j��~q�x�� ����3Ec1�w�\�r���&�����d��f6v;�<���^ai1����T�'��ԞB�������t��L5+Q����ccN�N1��\"�w�Ťӂwgq��W`��\כ�H�8���Ȇ!%�F؛�{�L������m���%96���+%�j�R�:ڛ�L��h�vN��piBP_��.�7��z1��g����E�ԫ9|GWh11�ְf��z��hŹ��`m!*��Ԡs�29@F�q���?C���3� �;���B�!��j�Ad�P5���7�E'<�8�߁#;��߿���-m�5{���u�uH���^��[-6�ɢʖ
}�����׮2k.g��g��$��0$�N����_��z�u:a�X�����_�	N�%]�wJ$�@/�um(E
��>|��u��)qE�rVZ �O�h��;:ӀJ�����9�5�$��Ҙ�����q��.=e.�Ȍr�b�%2���)�۱�vEC�F:�	{(}�������Nk*?rlӣ��H�Q/^`^y|)����M�Op�����w-��-�����ѤA>Ȇq_��Ȯ�ʯk�>�s�O�����/��+$����:~����A��oW�L�@	�v�&�h���ȪC�[*�x�S_<iTi�nA���'P��<5)�zpo��&iP���H��OR�/�;��.�����#�,%�Lՙ� ������ȉ���J�~dͤ��,Y$#�_��ۀ��h�7wlbt�P߸8�T跓W[����ڋ�Q���ES����wʕ���v�'�q�#~�NC��5D�e�D��H??�|�X>,DW�������1� �p�؞Vr�hS���g6U	�׋PO�lu�ey�D�e�ٹ�Ͷ���y7�S䩾�e���[eW�@�_��y����1��[��{�3aDi-�(��zVP�`%̒_�L",I�1��'
�Of$��pCۆ�E��d��R5�(�b�m:�4ȥ���ۻT��i�ҭ��ͯBrA8"]��9�Ý6���s~H̝�=��1����X,*�<�>��x����Mf��I��pR�K��a�$5�9�Q�p*��eт�+SG(��N=�Fxw̟n�QN� jnE}X�'����/Oc�,(X1`��H��|�MD�uDm��J$Lr����FŤ���ɡ��8���@O�]�2��5ޣ.j���<'+9��_��1Y@C襙�V��ı�13��5=��HGx]�f�
���~M��E2��9�!���ͦ�����;�����������/?����.�xTHْ�����_��No�/��w�xh������M}Oq��$%ߒM�PI�.�Y���Z��tӆ15��$�rGa�ڶa���|/\�X�n,>��$i�X_8��l'���q��2��/�4�)i�ᾱz� '܂���=3�c�����G�rH�g�8{� q����T[��h4s�;
L�}�)�T���u��
1������_��eȌPm��iD��>$�p�ǫ����QN�ǰ�Ԏ,�K�E��6��l��n��O��j:b�`���!H<L£������R��	[N�%DO<Z�����T�Y�BB?��J3��"�����V�NR���^�ІDs�z�wB&�q�eg<.�����������W�Iq;0���c���x�Y\BC���P�w,tB�0̜�����(,��������g��&�/yڈL��C��֢D����	�n�5)�9©v��Ȑ	W9���'��C�)�G�節��]v�6�{�V����&22f�"5m�LG=�H�.WxIc��1,2&�҇�������@C"��Ն;��Bƚ�A�[��uݕ���mu��2���a������clMYNsp�3��ϴ6�H�W 廯�*E���re�����
QSq~�ݢ��ӯ<���d%4 g?$L�a^b�=�7�|"]��/q�����q��\�_8uoRC��i���W�,(4� �<�	��ڒݯ��)�u���0/�Ĩi[�+f�g�X'����@��3<J�	e�<IVN*3�5����f����}a��|�e����%���� (��wWE>�;F��M�����>d���0�,���)�N��׷%��7��*�2���BA����8��i�sOۤ�:��_�hbu�ұQ�Xw>�ۥ�+�\��o+���/���(qB���5>JC_�������[#�=���
�-�c���XzD�(��DȖk�P��ب���/�倈�}L��Q6���i00g2e��g^�͊Ih�f́�`˽��z��.��מ��&�.�	�}�ˌS��s��q��%�ز����O_��5�0فї�z?k�W�|h�yK:�9�Qsˮb������a@8�E�:�{1�X�}�t�LUpW^�z,Ds�[���0$�Dm�A��qƞ+�i�hkR���Z�3'y���)����`�|a�(���h�����_��u�"�%Dw�Dp�Y�
�+=�o�]=)s�5��'n}
G��<9ڃ1��]�H3_�|������K�$ �sa�y�9��t�;��Ua�p�9������u?(��=5�>�ŕ��UH��@ei�Q2�52AIY$S^Z�U���$[-�i}�i��A'�7�W9>�9�z���BDݯϰ�*��8�r�H� �E_��"�b�s���G�i��) f�!�X��icꜩ���嵣���K����n��挴���(޵F�19��}�ϧ��t}��^&����#rn��d�z��/."�L�í�wX+�w!Ǫ�F��U�{$@z�Y�J�����M��V���������_��7�V�����NQ(��^�)a�G"����mL��`��2� �U���J=�j�����M[� ([>:�����o(�_��E�^fP];]��Y��E�_���hr� �'�
(&t{��X��uK�R���7m[��8P�ҷ5��!�\��c<�+�HS�,�v���+U)��O��?�yL~��>���?�=�N�;&����u�����?k�Ņ�A�����Kl�ݘC���Hӓ]|�Hzl9E����"��ƾ2�E���}4�[6�iՔNma�[��sl���,j��Q�TD�pcY,�ٵ�F\��Ӊ��&]�����B@;^���?v9��,��ȫ�LtҶ2�pB>zң�XK܍��Ə��ְ��<�$���������~�]�n��@0�Vq+�4zd,b!�� ��b�h�%�P|gH�.VE�i���<�=��*��ֵ�M� o��Mg�0��d�`u�D������n^�3Bvڻ�*�ؒ�uϒ#�X+�Ůk����o���m	c�3gg]���Ć����(�D���ieu�[����9k���X�E�S严�L�pՊ] ��X�#ŕ�Z�$p4�#^����Gm�Shz���D��������vd� ����~u�ǣr;7��񄯎��h�&�6'ŵ^��i"����֓p<�7��3�*���$����!�Zc�(��Z�S*�u,cGxL� M��r!���'��ϭUKT��d& ���=�}��Xחf�t@eH�N	���yEqo�+�Tc1`����������㬉KO��9z˖ ,���K��r��_���ˡ��^{8g�D����RQ�vQT���ڗ�,�?M������.��/����X�a$^*i���>T6(P�������_���~����y,��� I��ӌ�ꑿ�yg
��-�_̺$�0J��F���H���b��QO&�O�,����j�;��L_&V��Ri���Q��v�*�Yn�եp��a�8c�ŒY��aE��5T�ab\�	�v���7�b��ҁ)��)�n�K��s����r�à&2�+�4N�ɿ�Wf�ϰ��������^%�g����0������A�����%5��`4�`���h�;���{L�C;���;����8�����c��Jθ��뗬S?��\pd��փ]����a|q.��|Fʃ�g��p����=����:��l�:�{���{Xε��a��������w�gW��j�����w����kCQ��UQ�{�7��޹}�.(�NaӺ��8DWcqA�ˋ<kj&k��i�Y��sE��	��S�	>�#�[nfi���A.�d<B</O�} ��Bfh$c�ޡ����f���%��-���r�X#�� �n�G����'�rq��.�Mϭ���X�A`'��]21fz���)���w0��
)�e�/xV3����>$�. 4��?z���yD�:���#��'ȴ���e�R����v�+�r����ߵ�]�����{ʕ<�8�%���<�K �7C�\���痕��>	}p�<���٫�R)E% ��暋\jx���Ou����/M��*�aa�l�|I�	�u��S�/�X�����+�	��˦�� l3M��1��7��9�����A�=*�ث,��;�.��w��j��ˋ�a�/"��=���f�ד�$�V'��G��uY�'�|{�q�� xwi(J
v6?����h{׎!���N)��j�`�f�zn��?�������D]j��Z�M���(@%�7��������R�/H/y��.�� y}�r= ��r���݆\b������vp�ިR�Zի��m{�&th�D�&_�HuP<����ȏ��H��c�p��:[����|7���w����8�`�xQҮ���o%�`7�0�dM���M����ٗ���}/��-����ͮ��I�5{f���]��-�*��{���=JI��6B�0�D��>�3-,_�߉�O
(�l���{��j�tHm�SE�w��\��3ۦ��n��%������'U�B%�uh�G1��C���pŌ��M��@���J�+��p���Z��z� O���|���S$���̒��ވ�Ͳ4��P}&�b`�za��B��7|`���-6`���$f~:I4@�7� ����Zꦮ�&R�Y�ڸƲo��*�����z�j��걮Sj(q�l'����p֖�+p+���%�ɿjW2lj�3��Bp�����U�3;�x_�oX);�`�d0�Ǘ��k�EV�Qq�@ݘS.w (+4���T^��Ze���?'�X�(���L� !��ĉP�n'�kF�oo���A�Ő��H^�'�J�����ډ�X�~�2�[%��Ut9������K�w�ʷ��j6%���0ږ��&��y�,SF _��JΊo���y���ąu-�cL�W�.`�cQ��΢|ξ��Qfݼ�K�	=��0y����ޓۅ"����>��F��� ����s��"V���`N��C� ���0�@ET�=�?Կ��$"-�O��=���Y�]k���<�r��� �����=/�j��?(����%2�����g
��@���?� �i&�I��^{9E�rp]ì'R�O5t���(��d�M���K���2�P����Y�U!ҍd>-3�� ���Ti�54r�;�뫇3O!�7F�aJ
���3�ޣ`U�?�/QM,�nf�E�`K��^u�}�*��D��'z��C�E$鵶C������V�u���_V�!�E:q�U���_ӯy�@��y-��E��#􊴤W��̒`��F�5�p���<�&��~��V6	Q�7⮵�swK�5O+�ƻ�'�ǒ��	O�Y��y�v�d�\4�6��L� �f~G����un���/����s�&R+��B"�]���<;�������8��m��j���dE9g��EM����o��9�����4��#�������c?���3���Hn��B 2�r�x��� �iH�Z�e6n6Āz��;��|�̮>�Ф���c��n&f����n�6�ad�I1��!3���� 4��̒>T��_^Ta�*�PFӂ��bly�ʸ�俹J������P,fw�P�S�ς�Lr(�a�v,ݠ����c�v�i�����x��)�`�섬�5��)�5�yPG�O�<6�6�q6�'0�[������Y�5��Rzn�k��[���q��\L~�J22^ؒ���N�ړ�R|S��n9��˲&6~d@�E�j�&�?�i�n��J���;!L��i�,��sI�O ��">U�`Gc�)E�a�^h��k~@|��~�F� QJQ�j�u8\��TH�Hg��̙*^FW�|���ˮ���=%�<��}�t����T���:�)��V!�7�uI���î\!*Ȉ��0���k޽�M���C��;�R������g���&�YOy������!�4XejD
0y`��
�C�����G*b2�����drށ��{���b)���K��P����w,�ÌA@qG���AN�$���Q�47�&=�"���j�e����Rҕ9`��0������������wѻx�Y"nΏTw�U���W�|��b�����S0��c �N��ݺ2�ߋ��D�ك�3�S~TI��plgP&q/x���I�P�@�]פT�TgwC*?���b�_�)R�C�7�|A�h�hm+���Y��b� �H���΋�DZ�
���{Hf>q��~�=�v�Fh[Ȓ8��H[�^���O�_W�����5N��9�o�ÿ3�O����� m�D=ww��BZU>��em���}V��t��=
r|*��~�/4|��%-�}{�K�na�Z��qd���D�ʱ8��-���m���� ;����C9'��g9��|�5i�}���ES!T�4$UuF�$�(jlWR�D����!���y,Zs�������$%I��(%��ej�~���ŧ G^rC͸����yV�$��1��{�*��c��4޶����F���~'<A���H.�	�N��ӿA�^ٹ6b�v��3`ԊB ����J�.tC���뻇�,~�f)heG�rF}�C��wo&r��xd\��1�qW�a�!�M��Կ?���� ����{h�ϴ������Z�j��K!W��J�8�Q��V'���=�~ՌG�!�
��Q����3����e��[U��.#W���F�Y��v�����W=���i�wd�W)�a�Ҕ���эS�B�:��˪�)�rkp���I5����q ��ׄ^U]�]ܼ������80�9�Hn6Aל�q����%��� ��D�M���K��_B��տ������T&L��7��t���f�81�mP��*��n�wL�I�^���h۠(�5<�rMib��5�M%%��T��St��+"'�n��� �4D�[%�In����V!p沒��b�-�f�7����
'�a��x�L���3<�5$����O�E<���L���������}ő+>�� t���e�.d\���ҁr�+>K�PYn�`��K_�m�N.$����SD�R{��E�0�c#��Ո�����E=�����'�]/�-\q�c��""���̲I	�t�P��[������Sp]+�]|"���AN_��z� ��;N���s�m� ���}:�U�W( ��e�J��#����1ᶇF<��F̳��n�5p�o2J��+��jS���7����87�IG'ֽxg S�ɦ��b�cP �DP����}��dUE��՛{�䣺t�d�\�l5v�"�a�V�e�2y����=��,;k�����z]I�p�Ò�h�i�T��8W��:��-6�~#?��3�;�Xu[�k�]G���B����l�ȼI�2��n��z-�dl��R��ZvE&���J/��'��ޘHr���wהՏ�Vٹ}D��ٿ^:�B|Qr<'o�92�%�޸5�<�K��z$��{��T�e"���[���wG.X�JҠ/h���l�o�J��{��h	�C
Q[Wx�T�H-?�g�wK{	���"eB�zK�;�-D?�o�I⦞��Z	ec	��2�4{`���mƃ��&�T�>zmj?n��d%�b�G���'+�1Eb�j���D�M`-��Hh��q[��  ����������B��,��T�ɍ���o���Xj`�<�d��{�7�$����tɵu �xRW���\�g��	��qو&A
)�5��������}�(:+@��K`��u΍�l}��X��������w�h�8䌁v��C�mj���#�s����g���X��;���I�V0�hJM����f!�A#ꑝ�y�V�_*$5����i��5'�I���i����H��p�����f���{�UT��l����T��PN(�KX�u1k�0g�4�BS�du����>h�YW����,D�c1L�oC���s�.����#�S���`�|��wzGXz5$Y߳�p�Ey.���u���fɝ[�|uy�Yl}n.s�;u�s�<2�h�u}�G�,�/�����>K� ���ȅJI�|�I� ���c)i[�h��w><�9�N؝ڣ����q��d�����E����~�^��A���-d:�sI�kOȿ�3z�OeTY�]��I  �GA�G �PXm@�H�Ƴ��77RA��-�e�ژ�1�[8�f�K�8]_�&r��"��� ]��_#UL	9�-����mZ]s����ԐS�;` @ť�H͢[fñ�h�E�,[����V����S�)���+��}ȝn6��+W�Z�]i��i��V[K��h?�+����d���1y�m�?��s}�dy%<3a?�����۸񕳌M����C�Q�8^�I�
%���x�7�m�����c�O�/].s��M�>���>)��Q,��M�uԓ�����C�Am%��`׈����8��J툵+����	��'M�
���>P�Ө~d�{�^�ێ٬�&�ܰ\ I���H�y ����E�M��z�J�<�f�]p��t��\�����@���0պI=�����`�y��*�u�f7��Kt!���#޻������w�����=Jy�d�ȕV��G��Z�Zwl�#&}�¡��E}f�?NTo����fL���S��*�/%s�aXԩ>��6�T�/h���F5	����Z2�r֟�5��{*[�;Z_fp�5�^��֢������m"��L[&�롫�_�3Q�Rr��AE�U(��?�:���w�)����FiP'�@�(�"}����9|�K��=�"�r��[讚*��No��Q&x/�dg(��lu�EV��c��I��kR������x��u���f&-L䍭�vݑ�;Bz������`��~��<"����8J0\��b�o�V\�U�|]5*��ăo����OD����2��RQ� 5b��<�h)���rK���	��
 ����"p�l���G�%�ՠ|�����K�D83�B�Ķ>_J�?������Z���FA�a�d�Kn�@ae��O�r���D3�'Pn����c�IǶ��7�5/@�u;� ��D2=�0 �A���0]<� ۓթ`��O���A��~ɿ)�dYt;�e�1�"dd��(�b-��w,Q��+���`d�%HP�Td����2����r����
�d�2���i�S�so����>��d���<�Ai�0�8@8���k�q.'T;�6E��H�ƆG�Z�'��{bҁ|+(]ݖU	��>[�;�c�gM�r����z��������8G@����Im�j݆%XC	_Pt�'�ޢ����Ђ�3W���t���ds�a4��?^M�4ǁE���'~B�+9���T���Ǹ��j�`�ٺ�(?���֠Z̒�֐��c���7�Kp�����I7!�'��A4��v~d����u�Uw씢L��e��2�cv�?M'�E�b�6_Gwg����]�HY��V')V;%:b(��\�Y�dh(n�'c�K�+�:& �'a�@Z��č�KOF7��fg�kx��n�_��S�KlFG���̭��q�Q"2�!M�e�$�����%)/fI�Ӎ�9"��rr�܀�N]v#ųр�"�Iǂ�叏�}�A�i��ll�������SY
��-�x�>�lZޖE�P�(�l��|l��,p_aX��su5�D0f��^/�۳/	�����W�0�퓵=e�ѼWuxw���敹��]�U[�<��'wo~��ݓ��Z���=�J`�G�Oi$�>�ۉ����BJ'-�c������ʌc����� �A�8i�8��
v1Wt�֝_j�R�通�11a��{�8�#'12��t�$\i���/��a��}�0��9�� e� �W>�y�<P��.��7m|D�-s�$���K�m@��LX=�d��z���_��'�Ir��0��<��ٍ��S#c ��� AR�z������/�� n��(�*��:��'�;���J��r����g�� �*h�]�����FB	I�/l�ԑǤL�Cz�vg��=r'����n���{�48���'��:Ͽ6/@�O���l���E4�g�d��X<<j�@��IE�8+Xz�
n�a?��́�T�Ë���\v��9�ģ�Sw#&����'�$jY$$���|�/~C�` �R��� ��������A�fYb!�@��C��o�C,u�pW��G�	���I�J�嘒*K�@�����.(i��2]p�l���Z�ŕ�2�١%��~�S�0nd���[�pf�&>h���(��!KB#�]m%��a���{r�>HHȳ�j#h���&�&S#��J���,��?@��Í#��e�h��<��OΠ�8��a0���ՌrD')T�h}H��VzL:vj޼���m� �o���j_���@��j��2&6TӺ?;~�60����=a��kuӀg%�u�eU	%���ܳ/@�=i�Y��K��+�}{��g�E�n=�SvJJ�Jr��.�H�=H��z�.	�^�d����7����<��3�`'���r:����4�ǅ�o�mR2����J����
�5tP�iZ:�C��<���)�`J�u����^A׿�2AS��F�$VP��,GU!�ȫ�hZ[�`b���u�_n���n�
��g�#ʾI�)\��7����V��gO�hR�����t�]�Ľ}�0*���OJE,�-�$�Q�Ḿ�&���o�~h�E��J�U*��0�����:U�8�Q�Q�k�c��?�u�x��m�e��ո�<�Դ��"H~�G_^�ML�x�H��Z�O\wK�`��"S�'	:
���J����'׌
�!��~�W?h3�4��L0�����I�A�a.V��j�M�m�PGi�HKd����K�SE��K�V��&�V�ܘ������jѤ,C�X�M�O�,��#*<��/8�jh�4�a�p��  R��&a8,E�
ҿ�׵�oE��1�P�,>���2Z�v%<�w��y����[�B��{ `�,�^(�r_�:zJk���ERI;�;E%�G�{\#�v�M�k��h�P�-�A��m���Qv�Ho Z���;�ΜM-uH�'�I( �$�fF�b�%t�9�g�6��ԏȝ}��$�Am�s��+��)��QH��ѠVi�1E���*��:$Y�=�>����A3���C[Q���w�S1묔�0��3�Gl4�0��Vj#�bMGӛ��*�2�Y	<,E>�vx�WV���V@�֢��L��=0P|�_&�J(�˃�������۴���1���j���nRw�~z���P�dyU��E���M�'(�=��7z���x�<�/�.(��	�Ҧ�<�]/���ABԎ+�{�Z�����FZ�t��LD��1�j��%�{mqd��i�2��3�F�!�I7wU�T��Z��tKq1�K�%��X;@��_�ݮ��0�t�t��8��&���	���h+�����ړ#n-Ǥ�;#���c��Y�,�u�\c�5+V0ӌE�=���1r���Ћ��1�Jf�g���{Μs�%�V����]<�o"T\�́�� �"n��c/Ҍ�k�.m�L`+-�KI��:�ѻ��07I9��`-Hԭ�'{"�ܔ��HZ��� ,w�ƻ�9@63���/Y;v�ҏu��Y)��pS�.��X�<S��P4#*c�>��<A߹nE�e�M��$��0%mw)Q��P�a�xg��y�"��k)��=
qK���jHtb��}�����=��U=a��O�.���f��RY��_kz XW�n�c��_���N_ߩ���^ �ޢ��z�9g��XT@��=AK ��ս���[�8I�ъ��p���F��Cش��/�iaކ�(���n�2��"�-�"���U 0]PjF]��L��"j_�DY�9�$�;¿��ȳX�wh�z8U���UǢ�*7��-.nf9����N��{�ބ/��e?>��`Dq��q�t���#��c�� o�fn���䣎��n�x�>{p�P��1��z��jX��J��$�ޡu@�;�I����:�AJٹˋ5d�"��6��S�ƈD�Y�������+������aQ�3,1; �,�3pD*T��v�ک��+8V�=�-�Y��p"���9h���\�͝�u%��0����w�p�^����D���R`�!hϊ7B�x�(��T�3C}�7!U�A����y~��>�9�(*����̙�H;�)P��Z��*$�e���\�	�g�l��lj�<%�Q� |<o�dC@gS)�W�Rn��x��&�������;r-rヤ<m���՘�韴X	ܫ@z�;<�^���<��xc_���q�]�з|��C��:��+Yk
]J?��8ͱ7���L�y�q,�<�V�{��&	X8Lј�����I1\긌}M+W�����9 � 5�Y�b(Bp��tDnl�Z@8.��*�I	̉��N���yQ�𤣖VJ�h�+�V�
�W���k�9E��thP��)���H�L;}!��P](]�E'{��[�St�>�R�_��T�]c0�*�u�Wͱ`�2�8�͚6�[���\j��`�,����̮ϠK�z9��af�BU�E�!�JoxU&�50vT��rV�I�/!g�y&����0�|���Fcҩ�/�4�ߞ�'$����+�'�F�茦"5�J��3jc�SW')��� ƽ��������`]&r�&���Dt"�X�5�S�����4�o���D��H��V�*
�k+����h�Г��sk��yҬ!�eaF��v��!�
l��ȗa0x�f���d����M	p��G��iv�����'T�JUQ�7%n�1N�̯gY._v<ޥ��\#��<�i�(������~f*�7U��E@�C�������as_uK!��o¢H���l�K1!�si�-G��&�`}SRy�g�#1�|�(k�u������	t�9�JBZ���@�����U��s�v  ���Y�]�S;��j��'����K�B��Cj~�E�F&E�hB�k��7l��t3<?P��˦T��sŗ�����L!5���}|~\ԞNpΙ�Fe��ǉ�C?������c#��k�0����҈����ĳ���OP��*68�]t��uub~(�뤍o��9��ݷu^���a-����:{j�|�$!_AkQ�i9�B7�����$-g�|���K�Q�����D��������ġ�yɅ�h\mĪ��W�O� �E���R�M���u�Vp�=�ץzw2��t^�H��\�U��ǜ��&�0P�f !:O�;`1q�O��!fk�<|�M�~��NA��R�*K�QS���%�����֓��Q��5.�k�g�	�6�{z�l�s߽*�Uminm����U�Yv���Uy����]��c+�o�h�Q��/ULބh�t_���V�s^��H�,m����r�qȨޫ0��_����<��'nLz��.M����%�RyLQ7P���U��ټd6�|�b*-w\<������i�OV���i���fj\(�X��"�(w�a��$�"4_$r�K��W�@`�I�;97��dzd����b�R��`@?.~���Ld��Jn�����$J�74G^XP�lh�vj��д��ʹ��x�����]~Q����3�r�~;��Q�����g��w�~�ͪ&���O�mM3�����<{`��H�oI)��&��ˀ�ܻ�"l�i���Jfjv��/��[�!�̃�0��*ZG�Q	��/�p��QH$�#�����p�B%v��N2(ϯ���b�5��8�ǌv�V�6[
�D����L�d�9��P�rQ~�Kt�7�	�T�sK��"x�:oD1d����k[}��`��i��m�*i�IM#z�Qq"����&�)�F��N��m7����7��T��R�!h���� 2�^Q jg-y䇃�^g�{p�zׄ��*c3����o>�����[v � x�f�@�a�U��ОmoNJ��C�N��.:.wa~�h�ZԞ�ꐣL�m� ��X�+�cQ+��3h��!�5Bب�hk��=���D�`�3��4�X�i��6e��b�Hzr���v�J^Ը1�;�b�g*����w ��=Ҷ����ƷA1��1�*�\ym	x���{*��r������`r譽_gq$�U��9����V�5f�_ڶ(+W#��k����%!
_�A�}�����\��Ľ��=�&dxy�3�"��	����[�$.FV�-ܯՄ
�d�*�\���@Tm���e���>����F��D}�;L���i�[��`J7tn�	_G�5T��c2��3Ӝs������f\4Y��:����@}���X��7��e�˸Eh ��Y�q'̳Dh��S@8#�=}�K��n���}�-=%� 
�@B�=���#���V(T�Xz�Ẕ���ք����M){8�o�����d�<��f�
[�·H//��ՃL�,��Y����v�~�b�T�.�bs��aף$�Ӭw'&��a�:fv��	+�e���y+7�^'��������k�a&gM��m{e���݇,��V
��'rk��3K�;��3� zᐖ\5ߏ�wN�Q����7��ڎ��23���f�L���Z�a�����������8H�߆u�H�Y'�F[oɁ�_S�q�I�7f<���S���j�8�+��9�c��p���+ħz�
��"{߫4�U[��Q�%���t{��f3�w�2��g�>�XH�żݛ�&A��\�M��;���ދ�o����u	��{!���2/o�'f���i�˽\��]�F{E6t�cl�..�7U���s]�6Խ�$��٠
\ϼ��*��|sU�*鋚�N�1�BJz�_�����G��E�?3`ɰv�	VU�^c�V/����K���H_DM�?#�e�[rc_P���aĀDD�Dd�kș��)M``E^��2mo���	˳�pu�(?����`q�8%���a4?�G��֋�/���0�4׺`�w��X����Z@k�V�����촑g��|�w����)يj���Q)E��?u`N�
��-�&%
o�����Ć�F5��]��1��1�|2�d:��)��}��L;��w�@E�MС*�6��4���X�Ŵ��cV�,I���S���ӡγ���_፦7������r5���NS���P����:��+�&8K�!D����w3����$��s�u�J]�������3�Xb�~Ā,���f]f�=T��&ʋ�V��Xp'N/QV&��n!�6K���Y��i��ֽ��;q�j�l@4�(Kd6�@G� !�_��U8n_΀� �}�i�~�$���[��95����oϢ3qB��SO-��Yb�w�t�Y����ʑoV�rPL�V�ȕ�u��pyJU�b2� ���S�b�Mf�-=���1Z0jJ����7�O�\Xڙ(�$�'�4��~���7�� ���'f����=k���ξ+�W�b�G���ʐ�䋟�g�3~[-�4�=������Ku�T<t1�#NU�a��;:�T�$�s�m0kn�I�&+��Zg��:+'�yM�ܟ5Wi	�_y�o���z���P��gx5u�k���|D& ����~qؘE.���J.�jIF��׋ݭ�I���4\	%-�K>�~�
�b��2gՁ� 7_K����V�q�-J��/{���7�"���]
>���"eÛO#��;�#� ���ĉ,�&�����C�P��r�n�7����G�KˍN�?��	�������|{�A �S�
X^���$À�g��ߗ�R; ���[���$�f�g ���"x�4��V@K>)�#>%�׽VȜl�;��ך}������;��r���.��U�jA�����^�(�� E%t�׳wFhϊ�#�,x� \E�w���0��l����
��I���^�Z�y')�R^��q��m���a���R��|�mӚ8ʟ�Ix:��L�v���UV�B@MO��dx��^Q��GGH+y<<�s�q�����&FL�ԫ8��f�h����4��`[�T�%Pɭ��,}���e��EѢc��
xo�8�N9��m�ML�<f���ŉ�����?V�H��2m�7����f`X����l0�l�n�eqˋ�݇�b�F�����cX�P��Sfv�e����6*z��z��E��'B<+Ϋ>���-��ɸ�\��Akwl�8��+	Z���3P����~��^ޫ���~�e�r��x�V��Y���»T<�x���Pz P�$�x�b�� 	��<L���'${��Ä�>�R�<���F�u.�Y3� ��v�ZN�!B�G�ՆT	���/	V�Pn*p�Q�C�g�l2�g8����4�����%��Li�)�*�T�qZ��� ��o���#��j�����̭��,,�?�Q�ި�%}��A�U�-��ȝ��=�$�p���38�i���G�Hm!���:��	(��Ϭ�ɹ:�{*e����Y{E�t{��%�m[���$e�=XCxs��k_DB+���CIp�� ��FMM[4i�0���9i��l�(���$���A�_+↑�@W��)��~T��f���S`���h*cd�@�>��A)OѺ�C%�ʦ�V
��f���[�B�;��L��et��;dϷ�����A�L�]��^����V�7|�g�ք򈫺�R~SF�T�a̜���,~1u�;��:�H�o�)�s��I��JP�O?�2�m�	Ĥ�=RXh�m�Ž/�<fܟ������6�a-!	��M5�OM<�p�.iyk��6G}	n�*	{�����PH�c��A«EG�[0�@��$�Ԃ��a$��[�������=a<:�O~,��ӳuܧ�N�/�OFO���/�<������ں�;F�(�'X2޿�T����+��{|���
ܰ�Vͩ'W�Fw�� ��_��%�G}��v����Y�ڭ��wG��p>��AOS���lSB�'@E\�A���٤V�L������=�W�\1������>�@Xh/ϱ�$�9�4�u-�1Jjo��Y�	�]��Nٴ'����Ⲗ���]UL7���{Y,��o�2i�%d+"X�Y�_�PP@j�L��>b�^9�t5v�}{�@Z���w`�e�J�q<y��r�9�`ȗkq�ٓ�[�(�f����X�sp����3a�&�ܺ0w̅�)f~���R�
�%�I��{Hj�&��j�a
��T�f��8;�h��k��������CP}�9F� �h��SrJ�e;d��ߺ-�'՟�C�ʁ!=T��"����M���9�;���,�<,�%�û���g��h�WM����X,�VB��I����b,��c�O�"{K�R��d�!D�p ���%��L�/&{���C�+[O:0y2�`���9=X�v���`~ �k~O}%���=�'�|��?��F��y*��?����Y���e���d��S�R6r��U�J �գ�$)ࣆǍa�$9Lr"c�琚�4��2��hcjտ��0�м��hE��-�ŉ��޴�M�JԼ��/ASVH��R#��C[�K2��8�Ykէ��wä��d�Sݗ8S��y���q�OP7"މ&�A��c��8N�ք��L�AH�Պq�FRF�[�e��9��6�x�x����D����b�+?*���5����D�>ô������Jpg]k9�z��ӕܴ������p#��YvA�K=�B�	��I@3�+.�D�	�Ĥ���X6H>pz��D轣�������	�ۋ��;#'Ͳ��F�`��� �v��N��%��b`h�R�-gZGs���-�
��Q����r6�%�n�ܭ���;�U��F7y�����Q� ���%��m��]u�wk��� ��/C��-�JH���g:�1�y��@��c&	�OuTf��s1�����_�AY�����Z�~
p���-o��fUT��K|Z_ɗ�S��KA�K�� �?S�����}>~S����M'�9�8�LҀ^ѷ8�rJd}�Y�F��>��;+8h�88e�Ha0z]gB�|z������%�`���_~�n13��Ld�����xpٷ��88�k}R����>��s@D�Xٲ�jRJa�f�k����	&��]�JU3��V�h[�~6өbDA����0�rU������i����Fye������ds��<���P=�����.�d���x.!�+�i%�������[�s<��(�\�c#��� h��-��8�}�`�aM���\Ϟ�c<���ĘR�а�����Mk}:?�3V�T��:o��>ɉ~���B��gH�q[�3����3n���f*w�$�q|>����v}������S���`o�GɅ�6F�bd�AFz:���O�n��������X0�_���_kp���T5��s.��b琐���d�V'_}4�Zd���~�FA�gh:0$a�sn��
.r���>�h������p���/E֤#�+X�D?�{.VG���
XNh�wH�.�?�}f��44+�w�|���6�e�w�� ��/R�����)A)�6�q�Bk���P'��f��f|AF�$w�׷�����-)���9s^����v�{e�1:��C��1��?i���kjm��aFndA�Jf�*+z� �J%���4�~�\q9�S,��溞508�OBp�?�X���B {f���3����!��t[�tөI���r��|�����mz��*��!�u�����������	(QV��|bO�)�>l��_�9�7L_k/��|��a���P~ 5��A���9��+��Pn�D�̹V��������VZ4����P��7��ݤ,�(�c��oZ�R,F�l�9��u�Z����0�)%6}>�ҹ\�j	��f����� ��q��2�������^�Gyqz�ఈM|��ұ'�_ #��}��wܪyp �v-~��jZn.�h^�����&��X���q����c<�*Q�|��q�[�m7Lj��I�!���E�f�Ӑ>c&-���aԮ3�<Ρlҿ-�IPa�-����Ed=k���p��)̝����x��ˢ�%_���L��~A�ʣ�R�g�q^�o��g�R��Pћ7M���d��הƮ<U�-������=B-&�2Р���:z_�ו�!���]��x�w���5�і1ZA3�5��2*#�������hm�(�B��{��kD�v>~/k�)/��
�`+�2gRi� �:�_����a[ �g(��j*G-j���;�wy'�Ҭ�r��
��$}(�^3�}��R��l�������l�������!��""2\��b��������J�>ݦ��Y�8M���h�w��vSӣN���t�xP�!��)��r�h�0�L6wx�g�u�Q6^����I��F@K��sҦ�R�w��� |�Q��(�&	����[M�r����GNX�9�aE�r㎼����h�I��ͧdB8�V��b�P�ӫ�T�Kx�>t3;J���qV\A7���T4?9wM��{�p�K�XI���t�v8�&�
�.�W�Wx��\�_9���߬A���T��HN�R��ՕL���x���x���� �E��G���k]��#cO ǧ�VĻͫQޑ"����_��5�g�T�VJ�U��K�8�z��odc=�I�]Yh��M]���#�S�Avko+���.�+��t��ԍ7Q*;(��Ny(6��,��/���(��t#袙ͱ�i��%���6�;ׂa�	zͽ�����W�M������#c�=�ʮ��'~׬��;�Hf�+�n���-P�(]#ucd6?��G�Sv��?�G�����W��Ra��PE��:�R<ݭ���Z�>a�W��>3���+I/h?7��(��L�^��)��<�i�@��F�*	�v���߶�3s:��s{��v�%L1Q�ލ�]���(,�w�͢m
8�/�~����b���� �B���H�Ʉ�?1����{�e�f��%P���h��rn���Pt�&�TI��`�3��t���lq>�h�%ar�I�vaH=IO���?���ԥ'��)�h�lcC��f�V��U�h�;����ٯ�y���d��B6J�pP7­���ޏՖ�!e����E�0� W�LU� ��?~�Q�u�O�DP�{���?90h���G�ŀ���JU���wJgws��j#�-�78a^V���0ED�+�.b�0�ޛ�1��xm7�1�$������J�K�+����L�����x�b���O�;�+<vQ��Ha�"����GX_}pr��� �2 Wig��(���g��^s(\z)
��Z>��%x�ѫV0����@��J-�6�;��W���:����a\1[�|T�dʻq���Ya ��3�~���Hh�Ud�~~)�W؎"��`�8�1�i+W���ziH��%��q��3JS�{u�����������
�5��o����s3m�,�.��r*� �J�_��c���o#��W�Rv�+���7P
,��&�д_��5���9+��)������"S���U$6����T\�W�_�W];$d �� �՘�P�}�h�n��J�a�t�b��7���p'LX�Rr�m0>a#����"Y��VP�מ��Ke��ڼ}�i�Q��V�?��8�S�q1����ޡ��Q��;���2�U�g(�z:.t�}��щ�����	�
���h����m�B��wI��+$1 �D�������7����:�g��?i/Az�4��� k�H-�Y	q�j����u�3~%�E�������h�١/�@kB'��<C"b��0����Rvss��.��4���n�jNhpw�;��E��
��潀�HK���{t��RwT��%��ӆ���~�
����5�hВZp�5����FA�ʀ�X#«��ڣ;)�r��r�a���S,VV%���~��XM3gw����銉D�!�MD�s��v;o3�@�����
]�M$OQ���"P���`W2lC�/M"���fF�������D��R�&����ɉ�H��׽x�L���:eF;�8xB6x�^*�@������Rs�j^f#���<c�}x�8#�t����w8�������6d��y0�"��d�O�s�T4��:�m�y�
��~z�=�"S%�<�1��MV�@?ۃ�{�5
�ŝ��I5�4&rF���!�V�JeL�Y��x�� �M40�SzNb377��*aѸ��a&1���g�{������m"�[2��2e�C缶��f_g�7�C������L!x��u��(���W�I�٩�o�c��	V2�g'{2�����,�K�s�#i�����~�M�?d����[#��J	<EP�����v+�Yl�'�t�����Q֟�jYP�cd�������HҴ �8M���!2���ֻP���H�eX�΍LI]����_=KqP*E:$N�?��:ʲ����w[��rj�����w��<��x�	�����z��D���]��dQ~$�GS����pk���{�팂B��R"�ܠ?(*�TI�&d`n���&%��0�P5�(ǌ���!�;rJ�ʈ�O��[��IrO���,�~�-��I�\?���i>�ă,4�n��(2��(D���Ӿx%���8o5�zB��[3��^� ]Uu�6̟�����|�cRp�Ow����8����7���oC����xxO��<˗ab�J:M�H\�������|�i2ͣ�������佡�!����V}&���.}5V�K���A��w�y.���i�P"&���0�
!ƀ���ՍR����Gw�:��ZL�_�[٪A��f*�r�`l��\��� ]9��,o��� �8����w�j��5��X=.�c���u��$�.UT��U�۠?X�n|�-n�Jo���זmsd@2��>�YNf�O��ۈ�lqԡ9��x9��ͺ���pf�H䠧�Q�A��)����0��*�Û twۖ�84b�U]?��P��!�{�s'�c\I}@udm��8tfC����כ)�q�Xr"�I���A=�B+s����E��_��&ݸ����ft4h��*��{h�yHXt��9�-y�kn��Шw����?v��!���Oa�qƹJ����}�\`?͋|~��m4���(>�d�W����?��f�l���3����T<x�q#L߭テ���8��B��&��P�ؿ:����9�E��n��l�G1U!6��q��-ep��6/29@�Ɋ�'��#�t�X�J']�n?�qK>�Z�� ����x��Hi�E�0��(��zB��*9�4-Pr��WN��&��)�óT�JJJ�dpMs|���C�����ҵ4۳Q6��rSx��0|�$ m��1q��cZ͑����P����k\�}d�b�N9;�B��b�M7&�o0�,�F)�)]W�w�~kp-{6��b恴\��!P'�4����E ���T�	�*2���.T��/����p��b������ ���LD��5���Ť�<O���檡]�Swܬ�2@!&=hIA����R��*��NR��+�-�_�x�7W�e�ߟ��*���1�r�8b���; #�Q�'v�6	����\�b~��y�&_��%^�W~p����e�VX�?�x؈.����#r��D���[�P�e��g���M�#�1^�=�h�;������->�	�1 �_r&�M!I�ꝴ%y�(��>�7�� 4���'+��Ji)�t�ã
1,�n>�0��>)���+����Å��n�:~���k�ƛ�j��1��ӷD�?PPҸ�|_�j^�N�trM�cG���m��>!�ߧ>��/C8F?��~)���˛Cf�^��ĝp�7�r�P쿁������R�K�SDC��͏��w����2��S��|�=#���&,��.��D�A���䲙�`�F}p�Яq�}sz,�,���Q��3�ơ�}:��]OiG�`��}2S��CD t'~�?�j��|���m���4�!�4�J+��x��pc5$�'v��u
�Q8�nX��D� �3�R#/\�#��F�G��:����b��>�Ec0�-*��I,����5�Od�Hmv��BXg�g����'�)���i���ϡ��!c���\�1n���[|;���(1A��=�a�*TwH�!�66���zRk�3t�K�2�������Q�&���y���k�$MO7mz�?��sR=��Z�,�]��7?��v"������-�)L�Q�o=���r��y�<7���"�M\�r����h
{R�!�d2�W*	.�D�'�k2;�Hx��,����}f�v> oꜺ��8O�@i�-�z_a��<�?��~�.c���̾�Y���z<U�M��m��R�_4C3C�:6�d��~a*�d �C߰b��p>�-�������K$ݪ2�=le{'�xط��'�!�F���h����_�"�6�v�yg/ ���b�������Y�;%ږi�$�{k�q����q���l��/�5����؃�r����73}��c���'�s�H���Lwk�?�fr�w Xb�O�$[�}A0�O�5��.�o@�E���$��� �|��6���O��92�?���������g+Tr��K���x��X	s�A��U�ֱ.Xv�0A���6IS�~�1�����M��A:�#����>&��)��4�p����}��}o���<�p��m�bO�2�A2����3Q(TS�r����E�V�%�G!����:߼� ���B)�5��a t6���P[Gx gv9�V�n�-2d��6��Yi�X�KO��p��ח�(��Sq;O]��a��dK%�R ��ߤc+�=*�+feխ�G,�&B; ��P(��?���>��)e`#3c1����g�0sd��[WY�6S#N;k*L�T��.��f����eP���$�
��ۣ��+�O�_Rq6e���ρ�%[�����7w��*�����3,ֹ���a����>T,QI>G���Wx.�|��ër$�o&WŌqtמ4�#���MV0�[��n�Z[�uŔ���ׯ�q~A���_�i��ǹ�����T��z��-Qٙ��P@ ���,��aKy�NO��a<r��C�-�Ni1?��6�e���kQX[q`pw�~���۲#�8��B)*��M*����[�;']�gx]_]�)� "��$��M1�&���k`p��#4�6m\l����m�C%9Ќ6��B��#{���]V���Z��>�;Tz����lk�;�Pyg@��f	��@���݊;VKս�"'��O�G6�4#uٞ0>�<��>��j��o�����N�o��%6���!�Z3�#�2^+�z�=���A(3�Ǯ���̮����RJ��8��v�#)j8$�̦�&��.|���Ie��'��VC<Dq]�#i0�<�o|ُ'N�A��S��$w�I�y�ړo���[�o�2�!Q��>�|�l�o�:7Z|f?�pl�������P�}9�x�y�svi<T��L�T�sMQ��RA�A����뤦C�w�U����r
$�j�@���e|�_�k����&�����n�]��$��@��)�F|�a��;kt����C~��u$�t�3�����F��7zeB�O�9����R)�g�1?H�7<��A�ښ">a�s$�Y��F��;|P5gE&(^����~�����7�]���"��^����g��LA5'ג��MF���r׵�l.��\�{i�)m?�<;���5̇I�$���G��>�OT��*=��z�ˡ~8�������<]]v��軥�����6�������L�oU0���>�yC6��@<yԍ�"����$��q��~[��7�L�3X�wRZj-��-�{%D�2�Nb�c��y�w/k��߹az��xX�����_��wuF��X7�rZȣ���� �y�S�n8�3������A��ఈٍqOKͥ���-�3�|o�*dV��yI@�/��wL�5��yo�6���8��Y����J�YJ������C#_��j\m�B��9�K[�Sq�ρ�l���pM���_I���n�^�;�)F4*���h�;�z2 �{O�s���3+���q�#��K���J����e�������"�&l�aK�Q'E��	��djO]�:�	5و|�`V�E��}*����I6����x�.���]3'('���l�T�ّ���S/4�ya'�EH:F�����p^������9�7`պ;�k�13�������'n�CL�0�U���|�F'1������F�Tbj��)m@�w��O��zll�C��;M�+��%�ť6`�b��
rPdU6�;�.���uu��$���x�B�?9V�-�a�.�3T�%O�%c��m��*�L1>x������J����"�����˱��7�[J?����3_�udn�*��kS�-E�W,4��u�#K�Yq��3�M��}р�	 �3�M���bx3�]T�r+%,z���c��k�������Ύ��9^¯	ES�.} ��cʼqRiw��~M�2�ɹ��:9(�6���
D��=�˴�֪�� ��ⶻ���yjK�
^Hy���C�#��PV�p���6�Z3�;���ZVh�j�㨮[rs�,/ި�����&L�F�c�ȡ�I,b\�9���}r��C?W~̇~7��0��utңc!�ÛmV���Q���m�F�;n������Ye��넁y�ҡ��Q���n4A8 '	�ڧ1R1��}ǐã�ъ �v����ۉK�8�&�t�xy1oD���e�O�@k�'��dRk=����f$g�(&�ȕC~� ����3��	��
t�Q�';�r�2�|���}��_�"$���#��I����=�o���@Jo0l�.0\nQ���N����7�\�$���P�1 �HWޟ�9���x�m�$;o9�8,�2�D��zD�Hx]�u,�Y��InC�����|���-�6��+�0���}qA�|���(o������Ha����11�^Q/���EdmLu���SdKxA4�#FQH�K	c{olu�S٥ �p�����S�r1w/Ej	Ы�.�?��3�O�{4���@\�Qx�1� �)k�Q�0���F��xTJ���R8����lX�N���N�~L��z�X��Sچ`��w&*J�D<�eCf�ڥFh����+�k�{G��'���`�ɹ������u����ZI�X���J�y��öW��V���@�^�k����>��ߏ1`l�L��������p���� a!���ď4�.��d���[��Q:@2����TH���<0��E\2��'e ��R��M���3�]�J�K碖�4D|�m�M�ׅ�X4\��� F6�&OVZjP�؝z�Z�;��ԗ�s��S�����U�?#��d�55�����'��-Znc�H�U{Q�5�<�^���K�C�7Ac�X}�͕k|HD��+Ӣ�bTNTN�a�(:i+~�|����A=R��h���!&��	���C�'�e.����L.�4s�j��X���'Q1q�(��3N]6���2�[�f��hߒq��,z�D�)��ZO���a�5����nm�g���
o[���#��auL<�Vs-�ءgJ���~2v�𕅩l��!��|J�j��q�̋b�
���E�te<nC���)�Xp���#�aD�xN��C�8��p���v�	�=���l���ND@;�_����~gՠ |���+c�SV�$E���.׀���iQn<��#��K�<��?���H�臷	��1Mի�nA�~�d�~��Ԥp[Ae�5�S<���?Q�8��$۽�'�P?+Z%[�E�>�bb�"�z��;4�}�ʠuL/�.z��'�,�j5���[_>'�"c�^H+a2g��Y<B��1���rz�ާF�]��$B�e�6�*F�7C_�G~����yشū��Y�R)\�����	�i��Lj���C��i�Y����կ��� �"�=
}1�fr3 �^&s_�����o�jB,��#��^T�q��nǨ(�n)0�1)�r�����%a�W�\��p0�ƿ�\N����rf?�_\gF����k��3���7*�MKY����ht��UZa� x�p.G�auDCR���D�Y����V��h*|�V�f*�X��iq
N�.:ߜ"GuC0��~F'��Kp�$ 	����SwgrF�P�lv���d+��W0J@��?�����[n�P�-��K6�t�E���tE��}�(�.
cJ��h@�\#�efި��pF������&x� Y&��Fމ�{`��e�����&���
u2|���E+D�jXo�3-���
�=��Z�[_��I_t�h��w+��=<t�S|�J��r��9�1%�3rϜ�0B�^��h)v����U���6���e`ޒt>z�,�`ݜ'�u$���N	��͵�8�d� 29H���Z��$og��ф���K�7'|M����B���O��0 �)��FF����HEC4֔o
ҁ��2L4�/@.;VtTީb?�ݸ/�͐ �6V=X�B�IAkO�����k^jq�Q�S����Pu�<� 1�W�b�B0�Eei𸒗�4=�)�l��*�jf���3.g�_E�J�դ��H�`Gt�x/@��/�����5�� ��9��v����{�A3dr�|�誂u�O�����)�*�@����ͦ��ƪ�%0��x-4/܅3��}�eҵI�|�T��@���EQv��q4�>'�q�O��������Q���Oje*@ͼ�_����uZ�$���e������^.r"ڙ�4�A]��-~�
�z�;��@�}�VQh'3�[V��]��^����7᷆�fA�sW�_6e���VG2�i�rq�� �9DFF�%:.��5�߇�œ^�"�5�̪�%��=���ak��!?�+�BX�xT��y�g���NĄJ![�"����<�4ء(Z/$�,�s��xaʡ 	2RjB[^��=ݨ�ф�ۜ/��O��oS?��;�Q@7�A;}�5�
��c���H�17��ʯ�m&�^��B���@
��T�Ɨ۔��L�<?2p�%�i�*C}V$�I��"�3<B̰ъD3�M�߿�z�c(i�UT�pԅ�P�j̅I�X��?�H>qsf��1Wv��B����Mu�Ub��E#��IŚ&p��[�GR&}&� %i),�/<ߔ�'�':6=Օ���PM�Q�V���W��4�J)b �������v�@*��o(|���kP�+�YE I7Ik��Z�%�㌉��:��g��b)�\d�3��y���E~&��C�����;T-���Ĩ��!#R��g�?w��U�RB9�RqXX^kft�Hy^�u�"@nB�gfH�a���>���w{�h2��u� �\�-crM�V�����*�of�����z���ͱ���L�Z���+Y;� 1���B쁶�yp龵(�CM�<��N��N���}3qv���D�k�W!�pJ"jz��f��<�F;˰�C�r�8g���Sn?PwƑ٧^���$:'NHDO�C� �`9��JZ�����]�])B�'O�Lؑf;.�5�H�ùf�/>ǝ�X2�$<'�<�~����i3m�����R�<��D�b~�Sz�9l�XK�5� 6�K�|X�81�Ue�BM�V>�릶��FoQP�HT�r5ʚ��K��В�e�������W����B��;���yJ�� D|�̴$����0UD��Lƾ��X7����+*gls���0P�$��	J�'�������[��	�p����1�5B����x�2��rЭUD�W@\���%z���ߧ$�S�2��^'�4�p������.@ˣoS�$�1��6��5O69��u@�����D"��NL=Z��72͓B#�E �X�ô}5c��:��r�:�U\���ش��Ea�C,��J�t�0�M��gǼl��,��M���L������o���.�V��q1��o�b��X�_�E��4L����\�s����K ���ټM_�"f�f����;���58Ȕ�Z���.DX/��~ y&o`_����fuS�K�����:�T�r�wks <(�zk��[zP�	��a�i�/�X�X7����%��(5��\a]#�?AD��|`������%�
>.�M����^���s��H��o�B.����рT>f��&�&��'?�s�#ֱ�ʧ��@�T[?�1f��b��Q�j%����6��0>��k�3��p/��)3�<Y����,�����ߴA-�4�|���n|�����j�,�H����eE[D@1U8���L��" 6�C�4У����<��? �Z�&\� F�@���3.L�E�sc�]�8�_��8��`������ 舊E�z1�EW�;��|T}�#�Y�3�������gFTM�>=���~��[��I�{�`H���J�J�qMp��(�؟��i���6��t�}�Y�o?c���eN�n�&��� �k��E�	$� ��l�%��+�>4�ʒ��]�
K�J��x>�>�/�g��&ijV�q���;o�O@pX.��<�I�2vK?�t�T��0%�l����}�.�����uF�kQ����oI�~�gt&~[��v{������HǕ��3 Y�w�'�Q&��|&'���YY���ɴ`7�VٙB��5�`�A�7�p>.�����u�gG�{�vȝ�QN��%?Z�ZAEدf�D�)Z���ԵG���Z����tEEҖi��{�\s˹#׸:��c�? �g+�����R�y������w�Cڻڴ��n�9��R����m>�z�{}*�,����|�m��CG��qr�sK��:a���4��u#,�i=X�~��.��I�j:4&���L����9�@.���?�嘀���Ȉ�FM�kA�R���(�����c^5?V��jodx�x�1�Һ*Xo�^�\^?�Ϧ�a3}U8����1M�����Nw�2�?�,�^���d��W���~xbyL�qٷ�[�`R?FzmNKb��g:�2�词���͂*4ULt>�N?V�|�,�]�� �V�ꋼV�tcKV��2$d9Y�y�yֶSԉ����p���|t`�j���c(rI��d]��{��\"����5�ޮ���[I�D6jV�R��0Me�&�ZOt�j�LYȾ��N��o*�%��F��Z��EXh��I4,H��a���KD-��T[w�6�J��!<c�m�P,�7��Sњ���q2����X���2]� 0�B�S!�s��B�V��;p�d(�L��;VR`&L��4߲wФb����+Pl�c���������s��2r�)�ى��S��n�
8H����1���b����T~Ȋp��y��dl�WBV����$E�Peft�4���I�9����<�u��k���6 ,��P
M��5�l%�����|��h����6O/��cX�f���
�M��;�(ŝ;�)�y6�2���#��uhMD\��301IO�Yn�d��|/��Tc�Eap�a\�z�����U�T�"^���#��<��P f��X��#K����~A���W+���.�������p�GE�}閥�%���Ë�Q�Q�1����a��_���^4Y��)�c�G!J�{�Wے�M�~���/��<��w�PH��� �b�17՗�mTKEb��.�a�G�M��\_'�D�lW����<9���;����~�������a��[~����@�1\m�/Y�lW�RPh��M�8��d�l�����#�኿8���a��6��쾗����"�ϴ���oc��J��nVֹ�s͚k*@ɘ���#tc�N4��u�_���(�>�kd4��u�l�¡��z�`��tZs�)�F8�Ȇ�$:���+p,*�tm:�/)���!2sSDx'%���E$؞.��*�W�F��|�S���2qP��W�x�2x_Z��r��/�PS�m���A�P�i�gٙ(� ��<߆�3���͎�yq���Y	���ʊBl~Ӣ��u���=��Td�A� 5�o�܇m�yx�n�3oKs)V�BM.gjqD��ћc��MO�,~:��lԥ����T~���Ў_u��N'�?=��#^�u�}:��=�yN��\b �W��)��B�Ek�/���K��坕	�ݨ���-�n��X4U1}�����5,J?�<<�J"�s����>ޭ���������,}0
��Jа���,?n�� ���<��.�6OV6����9��W4��,�`F7���dh����Ϋ��-�ǹJ��|'Σ��x��R)-x�����t�D�k��v�Gm(�1=���GgT�d+v��Js�,@W�&0ø�.�ۈk˻�gT��&�h���#���sڠ���ޔ� .x����{���u�X#M��������W����J�?��.@�a]�p��撡o�[�]��	�]�
��`i#k��� ���<��.v���Oݢ矮R%��)��Yyvg�F����}?�UL�VƢ}��-\5�.�T
���X�eo3��e�`Ͳ�Ǌ2��U�	�,@㋯��u*p��ѿ�<|�j���򾄾G�r����Vs  ���X̝��n ��>�r^.߭��I+IY��32*gf���5�Gԋ"޷�vJeQu�O���5�������jg����ܰ;�|>��L腶��߿��:B��=6��i?�B-��3wn���iѝ��e�8i�ei������X�u���3Ѷ�`��@�f/y8��3�38!����`dל�>6WÑH�<�q���k����4�\�T��T���d҉��s:>@,����A�!��s]�RPUTϔ,5��^M4�lC�W$;)s�\K�l����Q����i����̗4���pNxB��M#v�}�woGs�{����Kͼ*í4�W�˳�xX�� �eؽW_�	;�#Y09�>�`�7��la��JMoe��*�,���xW��ѷ'�d<&�X�;N�-�as�5���L��Ek�M�J,�(���?��P��L&
�F�	o�z�߉1��  0rA���vly{Y�O;��jr�O��N���a��0�e\a�"��)�󊳏h����;����Cc%:zf�5!]�N܏)����<o+g���oM3�z;�-\
���gË鈜��7�-?Wu����o���Q
��n�-�����V����(�kY����e~mH}�1>C@S4,�)Lc�w�gM���Y�١���=b-�h��J����O�׊�.���=ZO��p��K0���X�0CG3�&���,Y�H�?�}Q1ޔm>��:D>-G�m:�Y Dx�^��o�8��N��_�5GDv!+b+�i�e=�z	�+} VB��>*�QE7an=5uA�������G�M��V�st��1��U[���L/6p�T�L5���V����	T� ĵ��o�Gt�5�9"r���P73:I�b~��מMv��UgĞ�0���!	C���t8��P��&5~�Q�>�©-V��C�OYe7�NxFo�S��G�K�E˶[^��04(��h/�����ACb���y�Ґ�W�}����D�p[�%�or��ӱ�_���m���=ۼğ�&�!\�DCO|�é���=�|�����JL/2�����I�&�Bݨ�� ������I��Us�,� U|}'�mQ��᯵�I@-�-w�$��h��=��>��J�*	��QZ]��OCx/_I;����"�Ap�F$W�0�f�a����y��k���f�t�Y�O��E.�I�%���f�N�\��j��V�"@�n֏��}";E�D�J~nz�V�d�i��A5�@���s@�Ɨ�3Uz;���˺��w~u��(æJ�w�D/1rR0V"W}�T���������9*��).��h��M���%�͘�(ɻY ���D{����G�vX>)��ܷ�*MW�Qd�/>
!!���r�`	l6*:�o�6�͔���C^K����D�mW�f����ۚ���	�م{���.Q.�Q�oژ��u����=|=e��y�{�����h��;���j�{d��V�s���,��xȴ#�D�ϝ���CG�t+z39͌�Z�6n��x;#o��\��Sl+�GmT�朣Ex'��ݧ!����ʲ6�_+�2DSVE�����5�{6-�]*���Fk�Y3���0�5mh�����י���o���9�iv#)C=�%C4��OL>��붛o��,c0j�/�A�>���
כ2��[͚Q�/a�'rq={)�ǰ5�$DH�/�&O9lԱ�t����d�,��_� ��C��������19�I���T��'	�(k��7���+Q���`<	xt��:���:�;!��#D\��D�`����n	����):\,*�~RD�a����x'�6q~źӈ�d$VFƈ����\w)҃&�L~���R����.�H-��N�Y��4�L8�[��Ln�/��̔FJ �B5C�7�_$8��ۯ�|��=�t���V�Ԍ�N��)��$�ND�'������^M=���ϴ�o�_�)-��B�E$����H=5�Xғ	��]O�v\�#h%�h���ڃ������v�N��Rv����V?YOe�7��D�8J���zo�j�|["s��)�X�����UWXVw�Bp%<7����4�"��^�UT���=��%��fesŰ�\1���N�G���ɮ�"z�e�?op17,���ڥì��!�ƚ9mv����B�G�ޔO��kc��H���K}�1�E���B�΢�� &�u���T#����c����67���P��涭�b����*Y�������TrMO�������c����OP�����Z��ׅɃ`��c٠��KD��U���E���������#��rYC������{�����"	s����D�͔���oÔ����F�Ю@���{!V^�
��Ҙ���+A���Y�\确ƍ�0�KA�SA#j�|�^�KB���x���kH�3��X��Br*V��S����aF�w��n3��[T #�U7xM���@l55��'ZgB�����y}vLT;w�&;a(��ff.c��~��a�����pkĽ����0Y��/�y2�R��e�n�ҝ e�Dng�Vf��E�;����u�[��nf;C�=��(��pt������[���1m�`���z�M��Y�v��6G5bW |+o~�4I\
�u��q���~��c0d(�K?����;G*)��.�|�ǜ �O�X��٨��$n��'���<%l��\̪��k���>.j�C~8g����+�$"���1鮲.{�x��l�Г�YOa���R���&;�(Z�@R\��J�	'�o��`S}0�#��):��1 �ҮΈ�Lw����7; �q8��%�n��΃���I��+E�����B�6�(x7��'�.�\-]ۦ�'�+ P�gHw�&ih��D�B�T�J�K����"����֮������2
����N	�t��'`�:�_jG冷ݯ�l�ed����wd�"��jwl83���C��Ω���b�s��Η�����ί���K��CIq�r=����m�E�47�V��?T��u�K�� ۩Es|�J���s��As��Zi��� I����D�݈��Hг���aB+X�E���\��V"(��$(0I�$�,��0x���.��y�G���J6����ػ����N�[k���ӟ�G�2�T�ri�Is�2��206bh�z���ٵ��G����"A4z?�*�@uq��e��
)0愅]��P��qL>`�6a4����!S����!v�[և�1�]Q��P�#a�>]��֯[�`7/�&�m	��	��!��Ǩś�̓sE��ơ@��[Dw��uY^��VA� �;H	�:^�쉙ʷ�yx��+��E`�L>�����; �'�S��3�\R�$�l?��l1�\~/���*�.����n��KwqT��i�ѕr_y���t�eК!r|���)�	�$^u ��T����R?ܠ�M����S���m�ĝW�-f:s%�a�y�`��M<\��`��螷f}f�����|*b����y!�[V埴E���I�չ�:�'b���g@�C<h�z&������uŕٓdy1�\m��.q)
��R̍��W|�KUɸR8H�����?���$d|�G��'-�ƹ�����P(�C/��m,����۶2�H�V��0E}��KY����&�����òjp�b���a��4�r�5e0}㶉=/vI/��J�jz�p�
���{O� (�e���X�o���:��S�T�>��5Y���-(�$KL��6$u���0U����S�V�4y��ގ��I��|h�@y���REK� ʧS�, :��r.�#C���=u�W)�-XN�CӗxX�{�3�ɤ�c(�N�y-�x,��T&�d=��Pa�=T���bۣ%�^j�S�h����@%D?#b7����8�ٗz�3�-gdڲf���]
)`p)ѹ:��$hn�\vDVvc�j@d�B�bD�� �d�eZ��F�F��X��-]J��:`���>��Fڑ�pYG��h�o�ɤX>h$�v�Q>-��Qi�>>u D���Ӑ+w?�ljED�G����ɔ��[���1�RLd���#�H
d�~ӄ-�<,�[� ��v6�OPJ�'���m�s�����q�mo`鍴L�̯�M��m5�X������Z�o�}���QHب)�Z��?3��[أ�iKU6A�L�j�U���CG�l_av��{�&r�} �=�5��͜C1@��}�-�K"m�8b���5�Ի��Po�{�O� @�j�P��e���2ZL�+���/�zf ��B���< ��_�&��Y��1g?M�l�T=�&:+7iไ�>��{��\�K�r��-)����s����k��5t����N��\Ц̠4Hk$c %��@i
��vo[DH��9�kc�îU������6��"����m��I�GW��0B�F!��Y��\��"cGp}[e�ȯ�������0SYA&+ur�H�8��K>����]��5����e�N#*g���35�P[Tk�܈j[BB�(�����6���pK8 �s�[��_�~�^�	������Y18��{�?�6t�c�A�����N�{��Y�N��oFp^�|�+y>;�GxF��c��O�yqD=e�=Y���I��O��}��)��(M�jꢗ�Vu3����ï���wf��2b�]����=+ț��9?`c �ۣ�l�gru����c�2	� ���MT�	!>�%Ή�K.��ѭ��+X�%㭜���3�e�����'��.n��b?.��0�;�J�v�G�E�сY�׭�ŀ(��Co���)��r:�}]�]�V��3Bw}���pp*�N��m2��{E�1�. �����7��;��_Z��"B �����K`���\顶!�f�,��j²����/K�G��A��
˂��z�_�Neؖu���zi��3�b������v[Y��0�'�yf?s�&��y�D0n�o�m�����E���9&b�Jv���fDj�]�0��8l��p�����Q~��D��0u�l���H�L��^[^ʋ���ϴ�m�B�r}�����������.��J7y��tYA�Ѓ��W292TSKx��e%�J���JB�$�n��a�+`����P^b�����VA���\�˝M���_��d�:���e�|����
_�`��B�{�D�O@��4�}�X�5��,F��H���;�<O��w��D\+*�Q�� �65O�W��C�qZ�Ƒ�_O�*�m$J������,qO��m�&C*�$#7|@2���E/y����N����"���7��Ҩ�"�kn�?
�}��;�9��B�D�����0���	ӭ��_�f�5
��z��E تq-Z�A9��D�ͺa���5�4j�n�B�|B����/����Ց^VE���H����*lv�i��0l򉬰bc�جo�F �	����K�3*}̫7Z
:����u�t���
���AH��Y�,���a �qW���w���hdCP���A^��oP�&�rKc�S�-t{��}�ʦ�ۓqo�_�?����0�e|���%7���4��x�w�Ax)b�:�x��-b�O�Ii���'P!����<L��:JF:Nװ��E��z1�S+^������0���{�m���Ƶ�`��CȄ����	ΗܱNL��O����k p�w�v[U�r�>��<����{Xb��9�@B��&�4���	�oZ�b>y����夂L�F�@��,I1ɛT+*l��f_ �������堃jy}e�K[��o���!3鷳�d�@���νr+n|�����,rqe?:*��}�*�ݶ
��M��٦K7��ۗp��Њ�(̏c�=2K��WPJ_x��\xϞ>נ�� 8x?X�w7�i���0��+��(OF������gS|׏Jz8ӏ�&��(�w �^v�>;J�����Hٖ�]z�}ZÎ ��l+���ȴ�w$s���"�9�i��3����,D}�(�rDd��rKQ�X��¼Pemy�a� Ǆ�gJ�#��h ���>~~��E,�m8�Ҷư,Hb��=]�	�E�v��b1�e�+ɫ@2rՑ�_��4��/L�S^g>�'S�-#)3U;��������G�%B���+�H<�DF_�c���e�B�T�:tՕb���1����]��OL���z9�p�j?�7�q��?��C�'C	�jj�m�q*��ܙ9o%v����>���w���%}��ܲ�!���6��?J|��B]̹7�D�驱΁��p:��4y_�1JQq1a��VC�V\�e��q�V�ݖ.㓁�qIgs��k��:��O$�T�`Ѳj;�x����5�<��v��M�:�)�	���9�%�ݡ�7��ơ��W�%��I�,4��;���g�#���6�4�A�Zͦ��Nd�"e�E��#�MO Plo���9�b��f.����L����K�Z�Z9�>����o8*B��ǥ���Wm��6�0��~=����B�e�u�I�W�
�qs#�WA�V1�v.�2�ܤW�J��z�e�<g��8�Ďa�.g�(�����6�O׷y͹Mn�I$����bh�<xV���L�������:���6��2*j�t ��,L0�ѠnC����&2��R��z��oNWz�����>�>d�{4�-�����cV�m�:M�Gܜ���t: 0?=���	�ƘW%�OE
�b�f��ډ��4Y�6�E]�w����;��n�'�s�߫�t��E3Y=c�o���]��
=���-�^�0�e-�U��qݰ�]MO'=�C�U1�
��a���u���������.�����q��ɀ2f�9i��� T�j����C��L��:�7?!��q������70���Ttrr�{]%��4#_�nc�y�Wb�%�����y�_�uw_�>�:`�I1�X�@0;F��]6~h�׺/N�if�>0�:�#W�v>W�ڣo����8��$��2P�g-R\e����[�4�׊�RE��	���(��2�к�<|8�g	)"�)�v1� ɞ=s^,��,�.Z嵹B74@��{���O�a�eh�pQYyS9�[��mhr�c�M���h�9�
x�^�u���l�W/����\-1�ższs��Kͥ�F%?
��)�Ψ��N�#�jWk��M��� (C�O	t^�� �p�*C�g1�b�)A3�뼂��y)B�܆d�#���uo�.y* �C Ml�20k)�q����5�La} <��Q�cYL���;���u��K�*C�����]*l�~q"�T͞�Ї�;�H&��d�Kk��)iB:���'��h��������q�,(�L��^�X��")@��"%΋*4��Ϡy}�K������j���pD���^��e��=gP�g�<���I�6va��(ni���@e�N���)��y�(�˥.N�n�[r�{�l֜��c��"�4�>]g�����WzZ��D�=�r=�x�n���N����������'��_1�o�V�2~�����펤WAp��ۍ�G[��GE�%25"U�����>�ŁCG��@�V�'R�
	k�����Q�"��:<w���hr}%��I�	1LZ���
h)3�x>�23y'׬����A,���P���1խ�q%R͡�H��&���VR}�Z��3��'fV��~�Q~U�3~�wK�[��{`{�WC�k��$D��k`�k1@����j! �Gsz�؉e���LP�̰!`������+�a�c�nQ!ΊCG��Z�)�k_2������ߏ�G�u��o����9��
)R-��P_%�5��Kߜ�$߳i�qĺ�]�`���u�k�ٜj�*zN�v^�����@Gh�ظ�%�m�Û�Rj5��\�Vl�WOH�0~Xꘓ⽵J�O���,��V�~c��	�Θ9_��-�B�zk�p�]\i�J�9��HW;�2��.;W�5�Hu	�[j}4��(\b^a�K�J��p���?�L�H60]6�P�D ���h�02p�ll���s$�:dkTɚg��$��~䣚��Χ$����<��jo����^�V{�j_k/z��|_��{u�����*�I%�/�Q�pgN�ť%x���jM�t}��@��<���_M~Si�a�@�A�z�vYЭo�ɂ�\�#\�:�#�o�+�O��{�&w��U�o<��8:J7r��[I~
�ŋ��%b�$j���T�'	�Y�.t�e����\�9J���x��G�k̹�hi|��=�H��S�蜀\X �������8-�*5���Y��`�w���,�
��W�d�.�4�\��ܛ"8Z��ر��;�)�����N>_Yn��)7���5���;�;f��s������p��&N�?��,�zf�e����q����O6�򝰌�o�kW>�HYm�����	`��)��"�P[��p� ��8�_J�P��U9!�z����� '�&��{?���=1������#$�X�*ң�^�Ql���rc'I�U]Ҽ)42��%)[�L�ą�Y����D�|�tk�L�i���0;��EH�c�G��%K|�t]H7z1�h٪;�L!�\��"5��w[��I�AKE���{�\0j����$�A�GD�O����D�]j,�t�{3��1�<n1c��n��`�h���="E�^�#$>��/�* L��.sɄ�V�D:l�l|\�[z��
������f.`�p��؂���������ί������Y�R��t�\���~���̀���i�Ƃz�l���Zv�6�L�!���{�˷uj��z!��a��3%�P�V~�*٬��������#}�%&��[7Wݽ97�����oL^]����X)3V8SX��M��s��G��]�Ī!FЗ��̭�D��۠�����b�!Q�,��B�����z�'�t*��3>��R:>���ŭ���P��;�c5q���խ�D���5�����<�F7mb��cF�)�#�S�n��d���Sb�r�M쮜=,�&Ȏ��]ߐ�0��X�dt®�f����h.�>Ѯ�Z�����d�ع���+���T��y��duf޷�ޜ��+�]�\'ez���n�?)<�|����gɕIZ��Z�$7)��L��P"�ε56�su�t�ph�"�#��{`��J��m�r���vr�y9T^7���e�1H��+ӭ}�L���Zn��CoXGH!��1X� ժ���:E���S��M{�ϗ!�iL��;��gK��:"�+%YD���V�$fx�Ն�@=�k��ƽU�,��f�KI���`��h\�|=�G�R/��l���r��h�CH�?{YE�Mfxe [���'�2q�\�e�:��n��S;gR)Lv4A5�Z�H�ͬ۹x{1�ב&�͖����:�i�CȐ<�v,�u��\���r�uT�u?[A���H7����oA�C��� �C��D4B��)�=���d�-�1�+���@�Lۻ#A�>�z�c����f�x�t�͆��)�pE�vWY[񥣁E(�d�o�Y1�u`
�:��+���b�P��*@����{խg�m�M��>�}j�M��� }'���2�u�G����m�����z�:4�ǥ��L��e3I�+SH��DӁ����֐V#��ē�����f�9�D)�vHF4XY6p��D���yct�VRUzhn�� SϴR��Y|��X�E���s 	��b+��@�?̽�em�'_�PB$9�S�;N�������v�1q/�a��,Pi©Ʌt]�&3.�:A�m��i( vth�,o��rs�l�U�fu�d%�^�l�|��7۾�������WpBG�2�~�L��6�ӱ����J�R �1h9�qDHz��(hP�(FJ~a)z�e֮��`�8=��Yt�(m�&z*�� �ؑ�?�V�?ǾQ��~�ڼN�Hu��hQy�$�s�~��{�w,7f2JK�U����iH�4d�Jn��`}�>d��Q��i��C7��\���b{�&���y�`o�C�ԩ�JXv��T�W��O�t�x%������["�l����G/n/��ic��77Źq�j�0��������4����I%%���.]#��V�q�]��V�Ma)�5A6��F\`eōfuli��,�@�F:p��3������gY{dd��f�B�M�-B�.+�~���<�Ͼ����~c����iT�J��1�8�W�������h�Ȅ����ds����Hɩ|PL_�['�˲W4c�8��ײM����_���~�w�h���ov:�&d���kvsy4n~�J+�B�嵶����J�7���!C-z/k3����J優��y��0%+2Q#�o�I�On$[v8���'ꙃtM���_Rv_W�w=]���qc��<�~�%��j\xNH@���p��)���J��@�í�ٟ��fԔ�f�g$!-��i�B�]G��hGV�ԭ����S���� =1C���B�^�곈�<Nc�'���ǲ�@���gq����U[1����i:�(t,���(ep���B���V[۷��D{nD�p���FZ����DO���S���Ң��j�=@���^',61�^��-D:�/יy�R�h`�d����� MȚ���.���?;�à��#m�5�x����v����W�ɲ�Oq��w1�ʛ��3t��������ދ~i*+��FFhBq�!����k�����m� �m�4��f89�뇜OL�D������x�IMH�ֲ��9��9K�hBD�-�L�:�\dj]n�k�G{(G��?����ob^K\�̟�C����x×�0s����m�1���Sz{O����qS,���4��&�������3@4{��&�(��7�������Ef	�7.�5���Y=�ގ%&�·��PE������B'������|� UA�Bm�>�z*� ֈ�4珘lvэ@t����w�w��f�n<�>�H��@�� �إagT��lh��h�l���<��V��eጌ7}F;�!��1s�Ll.���I���RF��� l*�N�GUY�3;=nbr��X�K""g��elFK�Q�$s��iUVn[��Y�y����Q�;	��2��|�Y �E�+��L:��������Yh�R�=�2X!x��l��.��>����L�&�UJ������H��B����� ȴ1���2����?k'@�mj�����m�k��؛Ww��,ޟ��C��;��E*֡/�l'B[�[��%���:b����9CǈX��{�A&�F\Dﰚ���7�8�fZ߲:��b��7�A}/
'�gu�H��B��j�\�&��q�m/����tҐ�#kB�C��%��1ĩ���ᲢH
Ϝ�	f Mτ�=���m�~�N�I��D����W�*����g%�rR֗����Z�W�I}�����4�F�@� ֞�ݹ��ކ��בpa����R�`�a@����\Y��8�@\���z1�P��`p\�zP����=?:φ�W�{Q�m,P�=��(Z�+���r"��N5��5���v� �e�)�Q1�g����}��O��oF�����]Z�A��ȋ2Rp��9hͧ��"�i���v!/X��EB﫠8QAY@�^���O�v��Cŋ�� �TB��9���;�� g�ԓ�@"���8�����Ͳɜ[�[����m��,�04���j���{�ܧ��,�:ʹ_�X�J7��^}k6ݒ�=��LR��늷���tS�
����.Gw������x>%�/����0�OS������+�8
*���Q:��]C�#g��d��
��b_�j���o��KD��`hxh^p�~xD�n;Dm F�s�FÎ�$�"jmA8R�e�K�_"d�7B�L�Pt</C��zk�3��E��k*����
��0JJ�^N��N�^�.�	�����MP�[=��Է y�Ȱ;����
����.�U�,�̴�j�u���,��M��k��N[���i#���o�$��蒩�3�h_9"��"�	r^!,�z�LOc�1�L`�4b�ׂ���*?Z���P>)���K�&~"�%(�:W�c��v��d�g�,Q��ĉ|�}Gj�E�}̏D����3�ϡ�x��"���ෝb��c��!F�dP.�>�)`>�%p��e�'�tG�R���f��>�]��+TS��b`�b@�_p�D�"��<.�O\�A�b�-`/wb�ذ�	��c�:�<�(u3���1�!�k�ץ�gq��沱�����X�]��x�zN�GW�B�;�u-֬+�?�N���5K��	�z� ��ި�E��uzf� 2OɄ����տ�8����J������n���(���A��26��G05�ˠ���}PT*�AI'VH{����ܰ��!�J.��1L�󌰨����.�Au��F5r�V�y�&�7�&��+A���^&�q��y�f��U�p�#�Jl�>�/��* w��W�4�g#	ox��`��p�`P U��醜3y(�cf+�P��vq��O�3����c ��jq���j�о��O�B;0���%����>g�+!��6J٥.&u/���x�ڂ�x~����pD)=�s4�
]��=F�=��H(���gr Bq�V�+���pNM�:ijݗ- �N�XN�?Et�9��k�&���l`Ƿ?�|?�q�C��䛴�� i�7�����3�0-A�nŋ��̏���iA�hD�+; ZEgl�W�~�,͜�gԲ�/O�:��)�St�W6��^،���g��c��ՠCϥa=f�4�+m�� �u�e]A�ɋ!��[����D(��Q�z�$3C�B�q���DЭv��rM�0a����	�aXŝT�!n�>)��v����0�"���O��P�-5<�+�d	�'n����˝�+�++�Tb�4�r�����ꘚ	��-tZ�}�Q�,�f��c�#ϧe_00O�>�1y�so(Zt;�.�JvM&d����]K��6�3�S�eX�;��A������뀭K��w�+_���}��P��b�AHݒگ�p��x)�c<$9�X�P��y�zJ�ƙ�k��ŕ�T`/�k�i�?4��6��ܪ<���m���<�X> 0��?Xݲ�tfN˅�=J�?�9����`��p�4:�h|��#To[�s�j���yy�����$���黝�	��UU���0Q��H[�X�����X���d�����>!e�� J^���GL���6�MW�W_B�aP�Ł��=�,o�$m���p�D�+h�a������c��v�֙��]?�uk�?7 z|ǐ-��_O��Sԇ�nGȚie{7��\����K�����B���&�}�J���)(T�Yբ����ZxT�l����̄	���LO5xH���s���4���hE�n�aï�� %�<����x m�v?�����r�֭큑����Ѿ᰾:���Z>"�jV1�l:�����/���ե��|�8����1��2>4V>/c�K�>s�eg9�8]ǟ� t"ЁD��:��tc���.V����w'���l�:�� n��.�n-=r��U	�Q&0ި��GM�?BY�`u=����̸��;z�8
���w;g[?���O���#�1��4��R���8sQ�A��}8��\��mFv��Ļ��]{����9oTF�����G2p�L�ı��5����-1��]=<?Үi�����~L?]>b�r{Y���̏�a|N���pj�v�Lݥ��uW5D�Ǐ}d��a�Y�O������ݶx"`�Ƚ}�1j�|��cѫ�\|Aoܤ݆�OV�1�q�!�;9���B�o)4�Ƨj�=��i�B����!���S�Bu��S+����R��!��R+��(c8*���ͨ�ʑ�D�5Y-��|S�ܦlR^���^Ou܋�5GP�T�W�c�)�ί���������cH�X�$������{:��mc���+b8o�Rme��{��|���'��m�ު��_x�A|�PO��ń$c���9���o�nB�ga�\�$;c��d�C��(��r�������yKՏ��d$�FL߄�ۭ�L��@m_3ĕVt@�fv�TT�+F�W-�Y����r�U��	�}��+�;-qzB���$���:�U��'� �4ϳ3}ܳ���+ ����ln;G�'�g����(��M��7E �&��� B�)�ܝԐ=8�\�aR��09`U�x!_a����<��X�S�k�΋/��5�����!`0��Y��W�7�*hVq��.oB�&�e�kA����3\�ʅEԺ&�)I��	�Y��+0��K�S�2���`�$*�D��e�34�X߾V�T6ȁ�Md1�ivS��11;�Mu��N�a�_YR�,�l���к��Ґf��M�h�Z;�"�A~���,�GJOt�����J�J޽G1ID!1��~�?���UiU��u$H}�����7:}��t־����Ѽ��d����� Bb�Iet��*Jȁ:噶��7/����O[���ѿ.�D�a�Xz���~�T+��ā�:���E��^٦3���G�|q���. qW�����`3ǟj��9���J���ɰ�55�J����c.��Ɠ�W�x&2M�s}oz�k��Fs�����)e9޵;��\�U�n�)�M� �u�zҀ�?s���fOM����͖
ݾ�@�7͡ �H=@A��%���r���_,��x���^&����hGy'~�|G��{{#��S�^��k���6'é���&�>4��Up�����p��X�h�qג�%�V���:�d�={����%������]'��ɮj���[Ē��,K� %��:_��=�X�[>��cvF�O�kFW�:�g����pXfT��ڑ,�R��v��WQۙi%G+�9&��6�r���'3ǲ�[�	U��'�2�n�X�yy8H�`�ͼ_�ތ]B�ͼ�=�m�c�'q��(��g�葜=	�,N�%�B��w*�H�?l��Bi�k�A�e��#1�',��Nu��^_���s�)~�I�p�O�e��d�a�B1���}cI���g�i R"7�l�o�@3p����'V�Ma���n��'w��ݔ�p{��Q���1U'���.;EL1��2��)N��4��*��)�bh6,�·�h�i����S��X%��?T����%췰kv�%�������#҄$�W��"�����_k%s�Ji?�$�@�PF��Ѫ����"C��kx�M�&���+b���8}�C�����������W	BjL�{��d�Ɋ$�`)��0a�oZ�$�u���{g�� #ٶ��r��&b��po�!/R�ٙ�]c�T��z�wm��9`]�2�k̋U&��C�-� �(��֫Q"c7O\�အ��_��!(!%.��p�fpE�p=g../����P�}~�Q�������/u7�1�y��u"�S��u�Uc��k�%a��MD��u��X�[�qB�rK�b � �tȓ���~�H�|���^�ȋ�I��>�A���G��(�42��Ko�݌�VIs|f"��zΏ��8�""�N6X*�+A�pdC�Bp" lB�;�?�,E���̥��Э�ƺIɝ"��j�n��Xʜ��D7����xj�TA\�&cֈ����� ������ �]�ui]�$-K�0�~p��3X�$;E�)���������K2�������o�E)�u����SJ�K�4mNE|9��_ۢ�d��B�{x;�a�wP��|��xag�2m�Ɲh�݂ߓ��bP��"@.�,o���J��"|��Z�M)y?g�����%@߇Rt�n�3��o`]��Z�V1��l\֩��*�d%B�&�aGUl��[�;��[̈� s�u�Q?���,��+1`��
!T& 8�0V�]�=4�S¾W�u%w����`,��	��­$@r�=��^������%�N	���ba
��ޝ�%��3��ҟ��
�~��G�L=���,[u����U��?���~]��&l�g�Ѿ�?���E�����$z+ZԘ	��xw��pS�޳���ȕy^Zb3	�0�yM�L/{k�v��"�x[�����pf����#���[�8pNեⶆ-�����f\QV������ٓ{�?�r�7s���%2��$\��z
߱�^.�D��9b���B���tיrH\La�|���O�@�j�-�tĸˣ&�zK{���6��.�g�gyc$͢S�eG\aY�3^�wW�8'��i,����:�A�р¯�T��� 1�Ly/ǲ�]���F�cX��2BO!������=� ��/��Y��\���A'Ѹ�DM_�M)�x�G�nZ��#�r��2�XI:�P2'���op��V�O�;�fy�U��/�y.�/iZ�����PMj�	�1�x;5�)1�u4/W{L���6�8��&�Ң��e��w��/�v䘫|���!�I�i��D/TZ�[-u\��_�#��)j����s�(!���ۥ�Jd��������#/2uS��X�?fΦI[����"��}��=24n��Q�^沥�iG�<?1�M
�떀נ*1X����1�1GE73|g!*j�P*>V�y��w��Sq^~��>l���N)Βf�5f�4��?-�4p{}H�*I3=�v�*|��%$ꤺ�RI�|X	�R��3(�|I7��OR��J��缏�N�'�F�v�0M�r�!����s}�1������=�vL'��K"{a��Ň�ԏ���@�D*��0��U��A������_/�EׇU3�/'=#��zQ��43��j99�f����-�)�A4�Hq�z�ein���N$��Ȑ���y��e݅$R���8e��`�-����A��
�!+q��`�����&
��!���Aw&�#�?����e%�=�?W�72�H�3��b��&Y`i��n��:Vy�����H�^�ީ[��B��e"Q����������������[���RE;�S-%�ܺ��e��Z/���j�uK�:�w I��Hj���v1P
�y
��L��n��(-��9*g�$?��. A�kU����.���Ќ��E�4z)<����!�&PQ/j`1��`-?�F#7���Rj�ۥ�cz�Ya��(g�3*X'�	��1+y��Cҹf@��$�s���JI�,�^��*X���
�`����b�-�����5���1s��j1���gH@'��NYI9	|V[M/�BS}�ygu5H��A���8��vŃ��G/��I�?�f��C�.��?�nw������[E�
��c�g�J����k��筼�|Y�Cm�}�A���.�O�/C��4�m�W �R�C�S��j�G����x����~�!�S^�|ķRD��X]��N�iH0�sg ��س��'%��I7�K�7��"���Ր�k�;ˎ������@*`ā����o:+F�$ޙE��`<���rCu����P��Hz7�x/��]v7 ����:��6_��k��3Ӕ�,��G���2^�.�;y����3�58�����Z`�>��/�ѳü m�lݿ R���ỹ4�/8�����F;�5<I'��ǌ�B��������\�g;��Uc���B��c��N*`A-"�]R素m�A�����qe�ʋ��� ��4��2qSn-�#�D(n"�����z��E�Y�gB�z�|w��%�F��K>t��m6�Ȉ�x���\1j��\��o��̅Ńb�Xk�)x�t���[v��d�g�1rg���yig�*i��޽�p�|��:�s$J�U��N�#aJl�j*{ɼ�m�ۤa�9�M��l?j��-��`���D��.E-V"E�3>��E�L9��=Q��Q2�(�%�a?;�1�$���� 9l�QR�����c�,�<Jj��8�M�+�ԏL,�H7!��[[�#D}c��⑔RÁ'��7]���],����`��h�z��@-�2��̮W!��M{�mG���R���j���3[KXM���(k_s/�F)�3!;�g{�p�j֏���B�f��Er��E�=on����+ɮ$�`e ���˧"��땡�6��~���E��-�T���	0���s��Q��K�/��2ccX%�
�(0N2��0!Y��_0����	H��o,E��!���q�O��!�{Ҹ7����O[h/CK�Ro.z����?��'�"�u�=�Ptst��>�<�p�~�}3v�Wk�a>l�^��s��=�v�sO�<1:����M����x5}��"��`���w�'��q�V�&Z�O˴ ��op�}>p���`"����Vnݑ�A5�J��Ғ3p����a���oV��|7qns�C0ܳ��߉�d��-��1X�y�߬��1�F#~d@-oc�)��_k}��b������&$��\�l�tIG�r�3�b�+��.�!���Ź-���� i�VN[?��F�'�U���3���V���\�ox��0�?�8��WU$©cb�h8N_n}�h%�U<���H�u� Z��o�7�z�^�I���Ҁ�Q�B ű����GI1Z��1�� ��ڌ�x\�����">Y>���R�^i�$�ӝ��t�+�<�H'
'>B�xй�9�ޝ�~��'h�����e.���>&mA��_���W�rB��Z��wt��P��T�n��勍��~�!���q�<p�mI�\=Gv́�c��5��������ݹF֠:_\��o�7�S)�D���
+<�j��x�����1rQ��nފo�t�C������c�������l.�?��{�J��諾���X��E�/=g��m�a�O�J���	�w�	�˾k3��������>72>�>�kb���~0~n��7���G���p��l�ޓ��ɨ[,	`5��N "R�)��.�|���+�T��)$Gl����P>{��_��/�=���L
�E���� ��adN�}d�с��V=���.��3SҦ�e��
���4�
�Q�ʅYH"���\�}�!�V�o��ea?M�?$�㗥�1�3C!�u;,��y�JzO��޽�j�d��$�$��5�Υ�o^�k������lc���ʱ�����$c4����1ڵ`�(N*0Ŀ_vrs����ogK���\�+�1�Ʌ��wD�Κ��GG�-�
8�܌��PL�8ZW���	DE������M�,^�=��!ܬΊ[9>#Q�{g�T|Џ}CɄ�^"�p$�IFM�7�(puu�j8ޥ$�r�>Gwќ�)�RZ���%�3�����4Ѥu�a����)M��^����8J�n�~i�卅ףR�n�-f��[\.w���L���:Yҵ�-n��N<�h��q��l��Y5�*�Lp��DⰎ�f٨'r���1s�?�曭}W�)�n���e�����ዛ�b�� ���F��L��"�9�H��Ҍ�`�3�y�=��#tU��%����
?�v��b��qNf�#�>��`��
�h�&�7x�P�E}�PU9:Nij�h&���9-�w������H��G#���1D��̔	]Ղ�T���A������5{��FR�w�u���K�<�.�g!�xy%<��o�z��YS#�W�z�~��剅��`|n'�K��]Aԓ:u���|d���3����ӄ3+��L���7i7[��%��/��s��NX̫C��@����!���*�H4p��<ِ�Jަ-�:c�%�f���-�s����Fقf_ł�yY�b9���zR8MLMW���	\/pw��{xL����I�� �� <��Dx����Q� ����
Q��}�&����uk�^�W��bF!�Q�/}X��}�����#	��&����Ť��9h�I�����wx�Tk-�r�[s��f�𦼠����=4a�x��Ĩbz��ޱJ���y4���y�~C�G�hC>�G wruSH�+s�(�-���}xe ucM\Z$_�6�a��o�R̆=;	<)*:K�%�z�T¿ ����+J^�Vu�m�Hr%;\����$z�m^���Ϧ<$&�"Id����^3U��0X�d�e8�\�f���8���;c͓�pD��{�IhZA�9P��
gW��������Q~Õ�\Z��S����`3�Jh���V9ӯtMLNYř<��T��E�F�j�n9�.ԥ7)�[��"9��=m�ޕ�����p6}?U�@��
8b��������T�\
�x��E�'*l��|�+��s�^�YH�	C�o5hC�Lr�\Uш�s�X7qHP`�R��w��TN|Y%���7��ɻ���F��謔�(�r=y@�\��yN�8��Zlۃ0���"ޔ#�"�	͊�.;�l!%p�L�ߵ-٢
C��:�PT�y�L�לoҀo� �h��"�����|��_�g�J���²�^�S۩~{��hR�Q ���>��}Rh$�Wa0J�\�p8M�:R>FW�/��"��p���NE��fD�M� ���:�:e���YU$�-N諸WJ����=�h���V;��i��q�L�qHG�@��.���l�-��(��1bwn���.�t���=�X�>���J��9KP4���!*Ǜ᷀":@L�+@��ۓ��MJ7qh-iM��عL�0˔���+8���P@7=������ ���0	:�t,M�È���#��A�;k��}r�|N�3s�s
��oyO�8�'2�K���Ւ���V ǆ�Y�)|E��,�j7SO���I�])��g�A~�+㞦 r��L�Pą��)��F�p֛��rе�#��e_W`:�WN�EgY�;�0�!dB�2%�A������eGܭ;\:Q"�ҹ�y�?�^5��ge6n��r)n)��#�s1�go�F��1�EQ%A(:���9�쿍āt�cX!,���L&!�_9�*Z���>g'8@h����h��|�p�
�}��u0[�#�MdO�0S�	�8D������a���� �Qx<�7f|{����`�}�u��/�)/�լ���neV�~���3l��7������'��g9�3�G�Ӯ�窥��ַS���Y=�2`nc(�dZ�,u`��ϒl�VJ��2>n�����l��������}��C��8A����
AJ�-p�#!"�9��#�+S�)�27c�	�&�����s��yH)�Ƿ���n7{�CVQk���Ťв�OK�������elo<��N���$���9�0��
�����J���*:;�4�4夕'�Ԅ�>R;z�i{yܶ�����xxnf]����5UR��͉��No��"��j�H;;�P���󶁊��}&��9N�����juٶ��q	�:c_���JZ��km>���ƌ�mk�-�ci)���p���K�f��ٳ�cܢ�e$��7ed���Ʈ|�yݓk|z��ܨ��	�ۤˏͺ�*�6���B0v�϶����@q�`�>��/���}�}L�� ��L ��P�
7�����9]��;vQ�b����6�K1ۥz�� �n�y�ԗ0ԏ3�@�@�qޤ�CS_qt?�S0�J����=��5'#��au�n�m2!Hz2iF����~w�y�  �a�4dLV��8\������/wkޓ>J�ŚoO����=IˠcF6�aL_[۪�s~nc:>�Po�*�j���z��ʭ�A���eVbt5�<����z'޾�$2Z��t*J���ҹ��.�W�� I������BY�O	؟�����GwJ�Ƈ��������UD�H�2�����35�U��t��>*Ee�h.A��
	$�z���1Fmg���R��2��͵[�`b��:��*㶳�
e��z*����������a[�����j7�`�	Տ����t8S�X5���^��-��`�� �mg_L�W��ougSJN���F�LC�b�N$�?l�A�T���fj����JVy���Rz�W�&����N��6~ց�*q�K79{��!.X���k�K�S� ,~�1{�Y,�z	x<���_�$Nq ;J<�X�LBLI�4Ĵw$�؞`J��N�6r
d�9Q ������c��>�5���#s5�!b�а��ڢ=��¶������U�1�fMac�U�nݻҠ�bMn'>��7k�J~��#&��R�*�b�ҷQ�7�\�F]pi%�'�U���Vki����=�,�7���!k�*��Q�Pw�r��E�i�w�.�� E�=q.����{&�_�A���6b�����!��[e�7���r��h7�
2�%�92�,+p#��ϻ7���:(��:��I�y�~�0�٤d���p$�n�bY��{��{��0�ȿ&�Ȃq����4_�T�pz�����ˀ�Y�0�^"��`�?��Y��\�oV�	�yɢH�Ɔ������X�*�v�/�޽�����b���z�i�5�=8!Ou��N�����6K�d�n=���4-�x��J/zc&��7���xè�����.E��S����+K���H��� �Xہ�X����SYd��aHf���9+jI�2��pu@W)Wk!�����!��(���M����P�k�I��L���o���Z�I����8��
�>{���Xݛ���AjM89 ��H��;?�Jl��Y��[������c�:5tA�6�r>�����UyAW��C>���l\�e�T�Ʒ�9����/anǘ��d�����E�
+Ɠ^�:n�ƖH��=9��Up�F��P�)�Z������YA����>���83�� 	�,$����L�����֨޹�sJr�c���#$�F�� \����O��E�B����4��P�a�`��
5/�){������jЭ�I2�|��{�z}'��B��nr��a�C`�jn�2E����4ӥt��J�K��}�x��SҊ���\�,\ٮF�HO�3�F�"h�Y�Jk��z_ў�j����R�c$l+��볕���YB^���D���l�!}'��x��dNEC����gd["���fBR5 �k���,'���8����)���+�l2�	b��������ʽX����"MAq�w���*�����2�ZPƨ��3+���Ѿ1�Zm�f�ܻ��o���g[n��l��D'��m�z�jO��>e�&�o7�/u�9f�'��ڑ��X�<���C��o���%����Ǉg�$��;(D�=˶��+�4DڤL(��k�C����kS*���ܹH��V�,�d�W�|��=ud���G�F�!ͪ��i4�[B��n��dX��FV�������b9#�$�_/�A����g(�I	��ȗ<ύ0p������/9�,qQM�V�h5�|G0�TiQ�VK@�r$��F�A�'�ڠ�bb���d��{�t!S���y?61-���+���L�&S%B21wIȱ,	ç=.L<��Y4_B�mm�� �貞)��`&��/2"��)|�ֱ��~1�3��d��?`�mhu�ã����shxM��)�ZS<�oݣ_)1V����8?.}��l�-�q� Nrty~��h�`�c!X|tN����t ������o\��f�}��#R�t��K=�����`C�μ���e�EM6�s�����*���>H��M�2U��^���ߟ;Q�.�?���~g��#��Az=��=�_���V�_��6q����[	���Iux>�m�È�K>_7�ɬB����n�L�ˊQ�U�b�T���l�
���a��)��Ɖ^
"�O���S;&H i(�����EG{�L����N�
o[�V�s�G����>} ���;!�Ro�m5K�6V����ntn� 6anCD?]��F �GҮ��N�!G���f�`�p��H�Z%ې��lD�О�tےYh*o�Md3.8�����/F���#�?����ʧ0@��/�y��J�Ѐ�Dk�=�.x��⸃󠆚��_��I����-LgHF���%�._Wd#��Ϟ����GfCA�ą������N햗yp\��o`���#ME�t��$2-2�{?��Ja,V�����#��wnV�E��MJ)��c�]HYêϕ��b�GɆ���S�+�s������p��#:},��y�����W!qj���X�3."��i{7 �B�16�-�-�,��T��(��֊�[=���]d'D�� ��U�KU�~���-�˙�K@G�ì��|T�R\a�!v��Q�Y��t��<�ܮ�f�+Y�3,o������F��)��X�h?��Z�|��L�>�^Wdq��*�:��V��=.�$��&!�f��a��$��MS��ĳ��&~H������t�@�5VG��-Bֹ ���.�5�7�,|e�&H+����"�>�(LX�.����ۧ���@I	�����zLG:�B�;U�h����S���g�R�)���!B��x�NgD����:#�(K�V�!}6Dx�c��2t���lm2kq6Op��ۃX�<�����=����J�%[݌�l�EI�٤�sf)�40��IT��aw���)����π�ׇI^�^����/��82��{߷���}�+��?�#���o��4]@���>�_��8�7���h�jj�ɒ��"zaZ{�z�?i��&��ԂI�nX)�cQl�B,�	�Gvg�G�\�A�.h�!0G���#���٦Q�=�\ 6��,ג�ħ��<b4�5�j������mHgJ	�x�vZ�b�9�9�9�1��o}y?���-����gJ��b(H�͈�Ǵ���z^�Ll�̫���v��k.���	�O�;������L�ֳ۠{���V�f�],�t������E*�V+ �Hhv<|��x9��,rB�&�r����lkK2MM�&��r�"�hT�q���u6�����ߊHS�k����+P{�ɫI�h��,���Զ�����U�Qwx�q$�[�籛5�5�������ت�[�'��5sx�-�����i��[�v�3��'��}�.y
���ts@/�5��@r��1�:��8a6xAJ��ǈm��hц�;AH��)~p"$7E�ۻ�Nt���TP,#}9dr�%�:��Wx� 1�a	GgkLb�N�	���Ru���U�G"�*Uф|g����:�O�0�eь`U�cs��N@�Yu�pҠO<*n�6�`B�|�ݝ���"�^C��W(�:�N�aQ:���ߤ��~#���{Ei���W����86_�����3�A˰]I,�n�%m(�॑D�/���rz%M�%Z}絫�2���e03��0����7�\�W��z��'9*�&�UGt�yf�*v�0���Yhk�>�/��+wj�G�H)�����aBw8Ep�Wtg���������^j[4hsIȟnN�����&bN�^мc�z�'4�6���;?
J;�Һ��6����B��N.z���d�1�V�O�D�����{��b�c�U:���?	cҋc�gZ�8�J������L�ϒ���q��c�f�~B�)�~xP,��dI&��9�A�p��5�fHe ��sd9m�	�Ҷl���}�URi�\�ݙ*qV�dL�7���-������M��	ד���bfR�_ekX��pg�b�������]J�����E��+4����&�X&����ɤk�k_y�OڙW���ƺ�<ε��	1�����	�XiC�i����X	8��@O���Yp�������V|���ސ}�U{Z�G~�E@/�}��\.0��bj�Ⱦ���	�cZ\�j�}��N�I�e��X'h0�� �7����p�ȗ)�@���'�*�2P�u3,��O��˙��C������R(��R�طfN��-P3���:.�渃�?�4��<�4���P҄h�#�$�'�o����X�G:���>�t����|TY��\X���O��+�{1��L.f�\�F�O8f�	09b[1����}&W�a%ffA� ?� �o�/�����z�Btn{pO����#�=|���9!v�Dm�J��/2�<��0��#�]�cx�m��h<gw�ͼ��'4�}�P�j���d��Lf��������ڌraj���$� ���M+�Guw.4JJG2�?a�Q���7Φ�%t�큡,�w���B<�L�W�a荰h��Qs��9�+��Y�W�d�YR��?P���퍄��m��})c@�D$�N$t�9L� 0���^�nK�V�{�"i�z�W/� �ش���:�Θ��ڃR�{�[��z��ܕ$N�,��s}|��b����4�y�gٌ���`;R�-j"��\��Ҙ<�?Btn�:��'���6P �O�X���xxk��4�O���qU�m�������Vq֐��2�ぃ����I͙h�0�7Ñ���f�]
N�� �+]�����f�ι(�B�ۦ� "��������yzZ�fw#�����v����iI��o��vz���e�s'$�I������`7�j5�-P��;��DgZ��a'��G΢D��t:իQ�%��x��Ȋ�V)|����&�%�^�|�����ET�-]v��l���rQ+殺��H�c�wT�� V�6$����P�@2���n��oiNv�D�r��ۖľx�[W�x˗�El��L�0ͪUUg���T~�IS�3����`���3I��[�9���f��ݕ%�0(�f~q=]
i@3b	�q�@ܖ��w+��U���.Ӱ:8A���[5a�A��:G���r���G�e��ѷ�p§�%�P�Z��r�̍S����=�9qW��o�f��cm����ф!�	=�;�MAN=d8G��Y.��*g�˃G8��*]V�g	0E9������|3�S��7~YЃ�{_��5#d�[hGh�\�q_�%6H��6Ep�&�D&m���y����GY�ӃU�sվ��v\������7t�Kf~�Jrii�����( ���.��lH�P#׽.���fSY�8P|9�C�Jh�P�#��ڹ�O"$�AR��n)r;ͽ��S��k�R3�e�m�D`�ظ]�8/g߁'wt�X�?:��5I���&��xp��a6��'x�}�H9�ݰ���ݮU&����{�����$T-9��A����h��q�mɜUԧ|��hu�/��0�Q$TLH�	n�l���05�/'|-�d�o��Ӹ������/a\2usj�h-ᴊS��c�.O��T�Mbmh B�#�@U�
�s�Ģ���RK�o���H\3ՁN���;�%=����n�D}]��U�.͔4Pw�B�F��γ=vH4�Ǹ�幽(�����D��"|��wI���r��J|?G��7�	�DVL)LF\�͋ �	�iu���kߠ���]�<���If��:�8պ�^�n��ĝVW��4�\�"O�z�r�!I�����$�6�Ȧ-y+�tv��<&mW��!<�g�f�{��� "ƣ���!�'S�>"�� /04�gLj4�"%�|�S������ V=��I�"�������
�%SY\�&�����yla�m����JFʪ1s��4٥V11�ʎ]��� c��ે��Jst��=�jƺZ����N�R��m�6_�v`��f1rܓQ~��J�:����#�F/(���TqA�_�l�n�? [n!nY7T�$�Qn��%f�ffe����n��,v)D@2�R��o=���L��6��}A4��K��H� ���Z�O��T�"�Z�fZ�5;*�/�C�/��:�g�tl���?M_E䉨��풘Ǝsdq�o��u�Ȩ��0A
3�`p*W��ց"r������hQ�e��:��m����e;t�R���i>W?۾ Z�D]ږ�����]d�3����e<T�6������*h|�ҕ ��(of��1�&�
#*�*�^W���s�6�d͖��_���pޕ�C��a��ߡ�`j?pg&{$��a�leQ�}���q=wq��p�w�<��M�a��as���VLH4(�Y�I��8�hJho��NB鹖�����4��T�f���Q���5(D71������""���Vͤ�b=�'��e��̸�R�yA>Ci��sʡ5!�n6h��?�	��d(y�4ݜ�)�iR���3�u)'�~[Wdn��$����>�ݳ	�V��mlm,��S������g/�:����C[~c�af�H��Z �H�=Z�i�Z�4h�0w����(�B�=6�OTy%s�GH4I��ݪ�1��pܑF�4��3��Xq��������3�n�1J:�^ƭZ݀l<#!��KmI;���ڠ֠]H}>�;���״�Q`_8�PC�+����Tz�{�E�N���j��,�Z:���Fp��WH)82B �yY��|n�wd;c �8��mL5�l����D�~'�Ʉ�(�G�p6�-�e�wIΛm����_ F���)8�FL���޾���6iPi��8e�[B�ke�4E����u��-�ƎU�A=����3'YY�e�W���G¹�k[S�6g�:��+�90�O���S�1���D��b޻�'��.7oί4Hrv����v��	ҹ*!��a�8�
�f����_�N�B�h�e4m�8!��cǽK��4i���9�> ��v�x��7�/Aл���T���� u�AV\�B���@(dAie����K�!<%����.���&��	'ϴ��?�=I:�(E�]�G3�Ǫ�]os��鑖Xp�%F3�<���$ d��A�F��;B��O+n�gܲ2˯�ƍ�Dѐ Ma��@Y�U�6���Jy�I8�c�Pw�+�yZ�����~�K�4���3/����Cށ���MGi�E۹���UZB��sw2��Դ���8����'n)�,���A� W��p# �7f�������\Q���<7�Y��)ZY���Q��V�P����/��P�F��4��.Ѿ���g��cP'��2|*w��R�&q�B��9������h&&/~�5p���f{n�@J�3��G�ں"R��}�kL)��]�6?�2-�nj,�a�����x6�w�XF,=�&�M���Ys�����y���$�uv��;F3�ڑ�����:S�Ċҽ=��q$�l�W��ުE��Mi̬%�u[\;����F���pJ×�{g�IdR�9�2Ma�/���s���{1q�uE����?��u*}���#�6|Lo�2��[��|�U\�;ۉ��a��1��;yDƿa�)���
4)�J�&O��a���qΌ�����&!�
�r���ZQ�8�	{v�ۑ�x�ǔ�գ&D��8�|)S�[Ӏu)}Z!��Ȟ���Q�[�s�M��C�/�D ��|U��FHp=���`Ҿ�T���l�l+]�Q�5ni]�9s��.K�0`+-r�,/�!k������ogd#Ԍ�kb�5��ϭM�m�왕������#�m9Q�W垟�S� ��9��,�~UN�Q����ETH��>I�d"���6�j"�gZ�>�s~��y�$�q(�K�>�?у��Z5w���h��]��X�f�;l�˫���e1�ӑP�N2�T����(n�8��l�Oj�V#f���:�_��.d}�a�j\;W�c��4��_�7=,+�hַ�O��p̷=sk�1��Zj�M�h17��� g��U3����-�Q����+/[4����$�M<��X<�Vb�����;K5�C������Xڢ���n��/;L����	�.���)�g���k��Կ!f�{
��+Ij{���0$�6X�u����.ǚ������Ԛϰ`�?�Ɖe�jk@����%����o��0����[U�������2:��/�
~T�`��� ���zV�uP��wG���t� FK�L�4����.W�,(L���R�x����v�l�����9s]���<U�/��/Շ�وfx`A�c�& k��j�����\uԝ<�%�����6"�mI����WY�0�p����ᐄ�:`�d��N�ą���k6�������+�#B� b5���PY�,��8�X?�=̭�R�u���o�d�(9�$�a���hy�
4i�v����wX�kN<[��i�p\Q£;� Xۏʪ��~E�[��:�MԚ��Ԡ�_k��n���ʼɮ����6�O����݅��$9�8�8�������I!�uz><�xGO,و(�"��Y����y����d�i�u,�Q��0�ξ'!�K)�4�8?I�T=_u��������|}ۨ�xxT��c�'0`�k.3]����Z�R��,w�9��&:�����K{�F�b�mn�8r�\G%	��Ebx�&-CW+�۠��}�]�H&�d��:!�ԏ��\����eV�C�!o�#�^'��n�esp.��+'���%�ܘi�U�"�:�W:a�G�x7������.��&�Ehp�������&�u#Ӣd��J:j��GW�Gɪ�8����>�<E�ca��FJ��ܼ Fb´D���W��Wwy5�F�P��#zz� ��/65�<�`�7����4�ȟ����a�::ۿ�C�;6���% �  :ld��8���ˉ��@x$n£�*�X�[�yN��k���S�\R(E�>��8�%��(�����J�<�9���mhLR��������)�+J�W5��).���4Հ� $t�xw˶��V{�9�h�Or��y�S)�&���_S恃�� �5+Oo"@��S�>�w/R�
Qkw����~���"�MH��G����R�#�JG�l�^�Z
���{�"��Jc�Ȗ�g��]�5ՃE T�.�DO'	��ͅ�}�eH�oɮ�� �������NOM���܌�1I�<?�� `+<�&Kt㔤=���M�l��n� 
^K���E��7�20pN�֚Z6Mw�.d� .fk��
�~�|b�J��SD�9�����:�K�hB�.��Kfv�T��}�1��@9���ZX^C+��	�f�#Z޲]nɱ��P8�D����i!�~!㱼Xy��隯lI1�Y��#�ͭX�r@%�9m���7�>��(�A�'n�[I`�Ү�.��vU�"��<���r��շ�2��"0����CC	���)�Т4?���dх��)r�p��#�w|"�b5"�a������b�m�Њ]X(�lJ )��W��_��E�����/�OZ��mV]� ��|�D����p�w����C/b�bL�_ێǉB�RcB8O���/����3��֞�7�^�_����?瞍'�S���e�3�L�K#���<i��E�jA�4� v��z~���1!�|���*��bM��6>�w�&
H:.��4ze���!t��g�g�|؀�[����g��gk;���'Ɛ�'fs���I7�PY&����/xw׫2y�
�&O7�@:�5Zs{0�i���}f׉��'��������T���(�1~kdI`���|��+1x|%�)��63h={8�%�ѡ��:�u���l�X��k��
�ۼ7�4#� `��i�[�;���:a��Og�Riժ��>/ �����b"0#��QǒJ,f����i���)\��G�_V3g&(N��_oU�O\���Xț`#z)p�A��(������!bV�<u�
B����CΪ�
o���r?��@�S5{ƗQ��Q�#S&�u��d�������E�K8k"!��B.$S1 \�OP���:�i]�8�'��t���nG#��R�(�; 3�<���ӓ5�4����[��f΂�O�g 8���@є��<y�9�\�9P���i~.:w�ׁ�TK�x�<���^f5��Êb��IŽz��>j.dT���"�� ���'e�L��d'�fR����6��+�$����3�K�������G~�������!��W'eWz�Hq>ԇHv��fc ڟ�O�5w�jg�b4�	��e�P~y��ԟ� [ъ����>C������Qy��4�qa-� �?nRb�nP=#c���5-�ӽ �t�*<�T�p;sś�U��/�k�"� kOG� ���Q�)T�Q&�;�\���pb$�C��@+��"���6C�[��Rdx4>M�Qp�p��-:(�h�<�b�_b����	6'2!(�\ag�KzФy��j�s�!U��Eǖ�d������7�Ɖ)Ep/�q[u������A�om���p��"AA�7�ڂ��nI�t����2�&��(]�^2Si�5U�t�x�39���v{���<Ɣ
���{���N�u�	w���e��(�=&�<��z4���P���[?���S��w�4G{��V�'���J����lp���	�zCrS��P���IѤ��WG}����u�I�	�.�9΂�ԔW	kyI�Q"k��op5��^�8�<���=�?B"s����zB\�ѵu��5q�Y��<���13�`2߃B�	�i{��75�˿��'؃'T�le��}@�D�l��@�U]?���[��[=�̑j3��t�q-#!�i��/$vqX�3�����b��,���t6�KMk8�ft-o}ZOR `������C��i
L�0���x����Dh��%�)���:� o8����E���Kd#sӜ�0FR���W�s�<6��/O踏�6<Ԓ��i��o�:��9�M�4qL�˻�D��؋mW����t�1ڒ�Ls5U���#B筄�i�Gw��A�[��^�A��Ӭ&wJ�1��*��<�p��f�dS'�M�P�������&����D^�#�/��u~\\N��-��K�~��Ƒ�2��C�Qc�]e�6�kB�ufBկ�-��< @=�}D~9��;a'����7���]�����=v �_�6W�X5�@b�Mk�6{j�&5������A��d��Y3��q/v�JG��ӕ� 2hb)8%419�˖{$j��r�*?��n���#�;�7�#XQo鐋��jIbu1�=����ںo�����4��lk{e2�
��`��Ǣ.�˂5r�ҫ���?n��?Q<�d�.q��5Q�,��ߌM�9��N�:�b
�l�ґ�� 2���\9������w�?ۀbh���,�<����b�NuLX�����PG��X�Pv��07'�BE�fO�6Qg�GD�K1� YN���_;Q�P�WǞ�mց�f����0�F�3��%��5�l0Ώ�-�۫x���mB��+��-��M݉���AG�y���&<&]ueٶM��:�q�}�`�q��;�~�n�ϨD�F׀���ò�*������N*�NJ��&�#nh9��GZ�o���D`s�9��|�|+�f�����S��y�3|�d���Z,�@�W�~kdCyLadr�+T�â��%�\7a��|Q��:�Rz+<ee�nyT�"�>��o�cI��d-�f?s��rb��_\_����C���I��PM�EP�J��8�w�@$�����F�h.�z\�5�^�&�׳p�Ƶ�M�?�8�o�_�1��uT�Y� ���f�a.� *�u�1�p���Xa��1�oUc��x��(�(�l�X������~��xأͿc�Ϫ�~������#���ë�N�a�Q�s�0z���iBǳ��ϕ�J�h��1��
"�5:��$�W�Ug-���]�%܌%��?��Fd��l��,U������*]?����b�$�/x��1M^&��hи�r�on[<�Z���{�e�l����9�BM�ųF2� �Np�ǧ�������3LMpN0$�2�rǋ�P�&M���}����ܤ6�WGKzH,����|�U㹶B�/����1f�;�Ԓ��dv��~�g�/���J5\�7�9���fe�W�7|�7�y��d���������y.����.g'��Ae���&mXҔ�����>!V�_�N�UU_5�e�����6�?zI) ��[:�d���ԟ�}�ʂ��b���K�I�{��I!�<������H)1;���̴��3�ǐ�)�9�\�I�n�Y�84�������E�z٬�ؔ��w��ߩ�6B��8�^�ڋ�9�#�x(`cW7w�X��E ��%+��8��y9\�0�}a	J\�B�w��HߏjT)pE��;+����K�B�Q����G���/���S�(��E��M�����<I����H�t���Sώ�_R�F��&�~�#�5�����,���tM����X�Ǣ�v\�%������F�;V�s��
�ĚJ=A����
��o��բe�r��ە�Cw��}�8<?u�6$(��������:���*^miE���Jg��0o��.f��B�8C@k����Z��Z�>i�b4�L����ŠQӀ���Y����q��"��bʕ*z/������P�H_]�P�L��d����K��8A��cu����r5a�AN�ZkK�\��I��f~��~5<����y� M>���������M)����G�i=&R�ǣ����ZU8�T�\M�@q{��H�������Q���?�Q���T\��y���1G}�� PE�وx��Lt�aX�>����P�6$^ɏ?�tĢ&�x�����6D�*���#���,�-�ڎ����C�:g�nXp���~� %���omM���Dt�~�D�ũ�U�5X�0f�>�8j�,�C���1\�叽s���?����wm]����>�\)���I50bY7!�=_�ZU!�;eJ�l?O���"s8#�B�C}��U��o�AfEy�ѐ减��D^k��+2�1ڂ�MZ%1�eł7����#�{��K�э�g�x
���I�B�8���� V�����?���U�����D�^�����8m�$y��e�H�Ix�	��F �+,��1g���n優����iҀ*�p����(w�Xa�����}���GD�D�I"K�mn
�N6\4֟d��Sܘ���T�R�����"qc���K-ľ�(%*�J8��ןDF��2&�s�ϧ��&��x��~�p��OE�f(>�q���Hޜ�L�}n�
R��S�>��u�3���֮ߦ���1�9�)���zh�*H���\�����鶄� p|��Վ]
���pP[C�R�ZL����i��U�P�M�͟���/Qȭ@3�t5��<T!1�V�+����g8-��G\uL���Y2|^�mM�#fk��LQ*�e/lhUS-�_w���_��l�O��{J���B2�6��U'u�1�>���q� ���+����\-���o����0�I��?��^|Q���� ��
�efc1���-	�;�c��j!��\���&v�
���m��A��m�ѝ��.�bs�|��2~���wl�K��sO�@f�Z��ǘ ���{��c��?����D���4?s�y�8�����]�\ŋ��Jgq��0��[N������8 ���;��d��}#)h��������8�{$^��B��g>���<�\�R��P5C��)|�t�J`[C$�,\ۈ���򍲭>�	oqg��j��M��mmC���"q���� /��)Z�Y��Vg}�cv)!�����99���+�J�r�a�e�n����i/�ͧ���~�K�?Bh.�qG����O��C=�֜ͪB�ӎx�1�W}1�3�K�6A�pv-l��fӨ�61�al`+-)�
p��4��n��5`A�f�� ��Np,SM�lZ�T��Ͻ{���j���(2]]�Tz��7����x�Rx��|`��^���-z�m�q���8f]����}V��{8��q������ղ6g������æ~��*��i�H
�ă���̑�@d����N�~2�&
#�Ц��g�)=�9a������� `1�����w\t�!+$ �W���@p�œ+��x��'��j�I,g�(v�"P�s��|j�?HN�
���-�c(U�*�:�@����s��/�0�-��.$­������ X��l��x��t��G��өZ��|�4�ζJ�'x��}�_g�뇫��>������H���1 �%��mLw9:d��N�6�Ya_�]��7E���pJ�(��{g���1�H�L@PRE"A�*&N�(o,�yV$z��ݶ�b�e�ljq�(�֗���?�OW ��;[��;h��{֌��i��f������a@�	�$e/��12G�`����2J�����rm�� ��|\�6�X�E� *?#K4��c@
Ť�.1�:,&e�y@(ָz�����s��7�oY+��@>�~�>��7����|��-�w@<��o
�� ��S�z!��r�y{^�Ud{y��~�����Q]8"�_T�$�}��@�6H��Y�_���n`��-�R�?H�Y��O[,5��q���<�rA��*�����$itgD0M���-n ��ҡu�Q%ΡZl�V�S,l
����j���E����7O��hq^@���sD(.��nӳb2/hmW0zZ��W?|5��+���cR$����c�+��0�dt�~#�����=���{�ց?cQ�a��!�1��g�|�9h��1]%اE=l#K��l��ץ=̪�~Uu�������S�C�y�d 4�s�q��)��~	�xJa0vY�i�)8�q�=��uk�s������X�T�M|F�<���<��)sgD������݅���8�%vo�-m�����k��6q����O��/�������)������F��Y�V��0,vg�B����'X��Ӭ��\�6�����wwI��@Ƙ����-I�kB�x�`!�r6�h���*.u���K,&����X�s������_��o$���qXz��K%!�3����!F6}�'�%C����o6HI�s}��˰�eoV��Н�I�`��\2[mm �{�/����6�G�P]J�Z��#	�4	�	�(��(M}Ȑ�u+e8��SR%Z�q&��5w�v�x�� ,��8�D%�_�H値�+L�nQ٣�+����ɥ��'�Vw�O���̞����C�8�6�b����������T����:��2��:�*�(�~�':��7w��UY,���5u�i�� ��}�P�Ч��+��Zu��C~�i��	�u�d[	��l؊m��\"�0����T���H)��M9E=��d��EP"s�����%6l%B[�b�9W�3{�8.o��|������&���j�ex%�^���W��[2�R'�"�B��z	��$�k^I�.�H���4��<��&��bZ�.VuvQ�X8��6��^��V�܂��Xc)�ة5o	MP�	5|R�O�s5�c��u���yu�#�y�S�m�oU'��Ѱ� �1�1��1�����０�G�(�S�����h���tn�c�~_B����)���m��e��X4�hI�y�7���/�E�ӭW:������h�_�����_��@����K�Q�&�g����/���JQ�A$��6� ���C|
o$���C��IN8�����#�r�2E_MhS�?T������.b'$7]� k�����A�D�l�~�ra_=��Ԇ��ir���Y
�HX ��>�CM��դM�uױu�_[�$���m>�.�[V"Zhu���;�g	���<H�; z�0����a,�v��L��3$mj��_0���ߌ�Vw�����/��+�3���$���zG����'��'�Yd1�sd�s�����%t-��k�7}�
86[O�F�fK��w�:�������,�����6�!W+�}Ԓ��D���v��O���qT4�[g���b|�F�2���H��K�����S���X��:/��L���$ƕ��gh6��!�٦��hܻ*�e�l_�C|G9�� ?�����ESj\���)E{��ѥ�"j�y{TLϯ1�z��o�MA�6�;}��r�w��vYB^�����A�o�}	F�^/�-7�Q��E���}�+aC�(����v�����Uӊ���a�%r_wɝ�v���V����'TK�6��{�yn�t���%$&�=�['�$bz�/i���[��I{s_�p�N�:QY�!���j�T�x=}��Я�)]���rў*��/CQ�&9�Y��C@K�LO� ʎc�����w&�;F4�v7R,�Z~~
����}C�'��r�)9��v&"X�E�����H�K�B�(X)��T.�GlB>N7U�F]�(:��Ãp�7� ��K���巛�ƀ�/jp-}���9��Wk��~�F,�u周T�<�qʇ1̓霢ϳN�Z��J�u�|� <B���q��P�²�ᜢ���U��%�]~�^2� �C���:H�6/�f��ì@�C~}�K�/n�������VX]�������ĿȒ�}�,�G��FϠis��N��O����<	�O�5�����Z������v�>Oj��h}0Y���<��IdUV�z��9��$к���U�~��e����E2C@�T���L�1�-�K+SG����*ntp�!�$3�=��4E��h��H�bj���ٝǶ�ҏ�2�b���`3s8�j� 3Ӭ
r �S>�D�̾N�����9-���V�?n������W���e6��ۨ]��U��6�@�5h*�K����3`NYG��J &S��ap�SY�7�����\4��0���;�c�ޅ'�/�.����L�<��4L�
��	����[o�J_����k�0ö����^�x0G�!��gtIQ�.;�����#��Ʀڎ#P�Cl�^�t�0H�o�1�<1V����(�W>�j&/q9l��q�f5�ßW��ʿ�7M~�q(�/�mH`Iu����óAB���('�4���.ū��	�;��ڻ��nT���2o*#�0۔��4ۚ��x�<��<p��{�~���R����Hu�T.
[1�%Ǖ �]@�����#{��ԅ�S�K�24�h�D=v��'jB0��6�웋G�_MTX�Z�!������e�?��P�Vz����}�	�yWHJ������q�>#m�Y�Yk�G�O�-=h�G��6��E)�]�m/�������ܬ��i�>w��5�5v��8����<\:�7�;ڽ�}������m|tą�.���/�^�_~Cn���s�ܗ9���o����<ڹ�١�y�-�5���B�q�[�q�p{�Ǆ�O����_���C�F�>����!(��-탟<6(1�v�����Y?X��~�aS�F�}ʫ��C�ٵaK��+�f#n�/ûKur�ΉB�[�P0+��W}+-v���ҡ�4dt�x�N-CqwB'>��E�f=�j�j��*�fօ��C1��~�����}NH�����U���Mh�)��@����S� #a;���G��#O��SdU@$(�{���g_�Sxaګ�r��X6�����7T�{�C�V���g����@��]Q��~,8�5����%��{��\�4��n��%��'�C�eO R�j^��Vk��v�-���J���������9�9k�0�p<Mu�j���U���B�8�K���9Q�Dt�z,�@��NM�ې+��Є�*��~�$&�(��Do+)���N��"~�u����|�:��}���N60$����tp�xY���%��7K';�Fi^zC����@zޣ��iD^����V�,�"����*"X�H<z�P��� UB)J
A�Y�<F.ɉH��iZ�0��5n$��*���
t&"��d�h�[�4�M������ghk��$$N$r������.W�9Hx ]�v� G����ݲm�N8����*6e�����#I����Y�^h��T��pٍ5%�%��0�#}UPw���u���q �9�$?Z#Odr8�&�I�r�R*)�r��۞ye��F#A�i���P@�'gul������"�`��sq�i�ʞ|�M�r�ΌX���k���	c����K'��B	'�o((���[X����п=�I��8}� ��,�k��W>X�}��d�n�z9���a���Ϧ��&d�+K@?O�oAF4`?�|�,�8p�*G{p������ܤ�Q��p�%6���@���y_\%�r8i]1�o#M��c�d/���!�sV̒+\��b5k�%�3���=I�!@�����VmC���P�����`|&�D�/��C�����,�@)�,��S*��.�/:�T���HXH\��Y�=X��$?�o�8��EXIn�_o��y�e
ˢq���f0n'G�I�,��+�&\����uL�+r���?��>��^�1�2�ɾWI�S(�Y �ݼq�,��;�ՐD��%�G|�Ki7��l�J�RC�ȇDkn���V5�Z!Lwk���ԄΆ���w�f�[�L^O�x����o~�H"D�ܣVt����d�7�׻��FЌ�������V���z��T������*3��D�\�Ux�?]�;&z5��"��,]��A ��D����ՆM�!ꋑ;��e���y:C��+~U������.F��99��ĪQ@���" *ť��6��N���q����a-�R}ך�h�g���ݿީ�����K\�u�,d:P���>���ƈ��%T�%����A%L��@ו])�� �(�!u�.	�ڻ� q���G�̚�������W��qY��}N~����u����R/[��.�U|Sܫ������١z
�2`9��Y�.��;Yk�6S��Қx�������T�4�>`m��-�koWsr��u� �B�'dNǏ;ע���]c�K�� �K��g�PD�9�C��c��h���������	����3��zl��E	�Ď�,m���A�[#�-��WI�ǁUa�o	2+�Y�L���=�T ����QO�&�KhU��c�����t�c��9Y��#�)�--*g�UF�i�a��	���t�L8iS¾�iva��CݹËI��ʡm֋1��J&P��GV��N���5]��;`ÿ�g܂�u���������L��/dե�na������s��k����5 
bz`�`z�	�>Z�����]�5@�����s�ӹd�Ӝ�E�,X{��m*-���j�⭯2�߇�QE��t�,�A��D�u� ��y3�.y�9�!�(��i��k�9s\AsSF�
�h��ΰ������DW�fT0����N�w��,�G��i*��3֤�,��l
=�.FZ;U��RIO���ֶ~[�J��R`�&xY>�?ы*+�=���D��bf��=@�B��.�h�J���9����u.���3�k��<��X-��)S���Ν�އg�?i���'�X���;��3Ԗr�]�Ԯ�2J�1.2�̏�&d�I@��j��T���1�9�RE�k^�δd�b������k%�w~���}N���������y�ؤy���������g1�t{��Z 7 I��}'4oDʇ.�MLD��Hy�� W C��O��a6�  ���Q��Ye�!DTځ�+���M3�`��ˤrWZI>���p�ta�.��lR�g��������	o�'x$b��F��=	\,Ee+љD�y�9�oa0b���0p6׿~��z@,���6��K����\���{@�ɒ�*ۨU ?נEM�sj����g�C�6�8sŏi�����N�>)��uNx��AN��},S���Z�����ߊZ��n�s�_����d�,�â#���^���[f���L�)	�/�EU�������S�֟�'��/���.�~�*9�/������X��d�=60� �w�N{�l�����6AL��[|���귱E��%�����e�6\PX��l&��UG��1t�!]����e8m��st����!���ި��YN�+=�ZWa?0����VE0ԯ*"�csH<��-��o!@3�C�9&ˉ�Z۠�e=�V%�n�L��@*n���(-�bI�u	q�,f)&���2�^@�w�,|��~�2�p.Y[l��n���L86�E{VR��LX�QLIE/�oㆷ�SfV�D�o�{��͆��UZ�轀�o���i�IG&-,��9+���/��tA�a	.a��/�Cx�Nm�&k��B��վrA����k��aM��h|R�{�8��&��gѾW����~�9��z�Xg�^�w�-<AE�x�M�tt��ͤ�#���˻p��?����_��4أ�s#�m�WBw3�晵�����2�Ϣ�o��/���/]���'gt���h�r����;�ȹ�����E�ws��<�@�|h���_�>�eyA1���e��am�i�u�e>I�e&`;xYJٯ�ѦPx�x9��@�7N�p��0�������2�&���I�A��P��W�*�f��u���2���B�Q6>��c������Y�����v�Y��A�]|"5�$aDc�;��Rs�gb}h/1�5T�	P�G�1�d�z�V���g����N=q �;��M����fnPZo�` X@�����\����˖L�4l���ǱK��{�p�M�\��K�H1�"f�����;��l:�6��M�Lmr?� �(c������D�|��Cԗ�tq�\�W�8s�,��*� �Ј���>�����f�}F�۴,���+-�������g��֐�x�P:��Q;F�$"^���S�Tu:���4qu����l�3�j����A('�T9"|d����ض��	c���!����a��!��2�_��9�+����)�V����m�«FZ��"X£G	������y��M�������;��a?�Y}�Ơʘ�PZF��V�`��3�G��E�e��xO=	�?�*z�T]s�w��� 7lcl�a���\$z	�yږNܜ�ӱ�y�8��)����G;ca=2��?]��VJ�-h8N�L��7�Ld��?EJ�Ą���-�@b:�n��Z�rM6f�-|�5?�i��F�JE7�0��%|E�Un��.�7�v
�k�q��w�-L2�Fs� �~P��T{�T^/�����K;��|���8"�ʨ��;����5�����h�N�y�j�P�����ۇ�ϱd|m�Im^�YN���ժL�cw�JT�,�k6�=O�W�	�lGI{s4{&<E`��aI���� ���,L��ZV��Ab�O�>.p�&���P�[�L��'��3��4���g,&9��A�����CO=��j�Д�kF���T}-i[ ���1x�݊��s��)e�d��9���qUx���&�s#�^���k9\sR�8�����j��0�9�^J����6A6���	$�����(!� 5{���g��M������qs�2'?;�O�B�%��pᔒ3�o(Un�}��{$�OV&��g�/�3scxX�/��P)��X����+"�N}.�t����N �A�i��Eֆǿ�"�8�C��oՓE�v}���PJ��)�q-� (夐�k{wf`d�k�3�� �^'�-xߐ8n�Ԑg/�*<=�67�`�!���'���D��!�P���9-+Ҳ����LWc��њ�ɐ|�I��w�xZ�H���PxsE?�Bav�&�|�ND���'���{�v%L#
R�R��M'Q��>��y" ��4@��~ʁ��Iu�F��C�bY%	g��y�,�3~R�suhy��{UI�6�l��u�߉��f�.�$#a"=I����>^������x#���{,G��tCG�3/#m��_�>�1��7�r+q��KH­.�ҹ���Վ�T��(�>�D~-؄Cr�k,�?`��|��:y����s�c�[_#���.�^/���z����rts��T a�
��̸���TcV
)�T�� 'Q�C�Jf 	��Z�a�{1f�XVZ����1� ����eH���CJ��HE�9���C��}Xvy,-���"~��2舋���EM��
<�y)~������E%�Jճ�<�������!φn.
|l�����m"���x/�הu������v�����y^�ڄ��b�l�$l�*w���gdȽGdG��
���Y#!�B������l�E}UÐO����m��nԋ`O�p��qw�0��x��6�P|�Ɯ�Zs�!�D��`~��y�����Iʇ�>Wy��<EʷeG�&�D�d�3�Ѹ&<̾�^o�ol� �/
;;[خ ��2n�`��Б�m�>���ِ�
/��YMl_��9�g $>�G����B{mcq��{��h��.�ˑ>*{�%�9م�d �:���F�|��Ba���Ψ�4��},z]\3_	�,�& ����	�礈0�+2����"���Z�R�U	�?xL�X�4E4ϥ���w֡�B�-$�]q����
袿�
��K�xѱ��D��Ǹ;2<��a�q���%�!6�L���ΘJ?������3�����׊s�b2���={�q��W����	d�{�j�st~�K�9�5�RD���2yZ����K�!6�������U�+�˗�_q�a.J�9���sY�
l�(��?�m�1F��ڮ�f����a��{��EǦ;�$��{c`D����r����	[g��UkҰj��W�"]�<a^����w����^�`���N
Wƒ$lٰ�l#�ĕ3�QW抓������䪮�����Ke���C�d�F��`F��f��睢'M�hy��4���^*���=�_M�)i��?�r3��b3����x1����Xg���������1%Ն>l೚86f�O�N��g	J`�'{l��}��`&�pF�:�qS��dTd�o���Ġ��h�BsD2I��@��ۼ��T����g7(%-F�v��wmc��]i�n_V��O@q�iω�����+��.�{8`w5�ёq S:֕�ɌHLk���f
���y}�����L�A��QX6��*:�_n��>|T��ү��5=B�%�Wn���N �E�խՉ����K'�A����<x1ῦ��
\4��ʸ��LS��X�$�ԏ����=�	�%���Lc5�7<���@�<�7zxe�Y����ly�����᾵���ئ�z��pv^�����������tɱ6P���E���-@f��� �!d�L:_���6"Lَ0+�C�� 2�|[6�w�Q��I<�6A��	��h~�k���î�.�+�,I�1�Wl���V� �s4|zĂ��^�Au!�F z��Y�/n�\]�s��D�����C�#R5�4Ư�f��/YޘQ�P���	�_�b  �Wr���_ꢬ+�GKZe�Bx�����Ԅ`���'��D�AO/ݎ<��8���O"�^�Y9&�⣟���m�R�l}re9�(�(ɶ�0�����%�MC4ʪ����M<�b�� 7�����s�c�K�Is��Ǯ�J�����������֥���G��p����Z5"P+ȬF i[�ˏ�xR��+X�Z�S-�4�K�g��Z-��h�!�w��D󾡍� �	Q!�S'-a����ę��p�=��9�0ű\gu��7��+6��;�}?�R����c�~�T����8B���[7���6i�2H��%ل���-G��v�c|.��Р^4��l	ԫ�
� �|�&���dʜO.^i3�F K"������'ǜY%P��`��5�ڍ@��s���fP��j�
0mmv�"[�#[�1�*G}B�ԅ�� �N�%~)���6
_-oYH����2�#> �%��2:eIK����� �EG%V[�
��k�Y��,�Qy&����4+73K��Wt��;�J�}^myé,�0*�r߂�1\3l�x�Ͽ����p���^#��$�M ҼT�bBL�����3m?$�<"�~�b*0��WC�'q��2�(|��oHu�Y�s����1�2e�ڍ-�0Kild�`���>�}���Q!sT츖Kܡ��#�%a��#-�!^b�;Cbgkc���O�Ѐ����Cm�V��&V�*a�һ2�.��-h{�O�fB]�̧�%�:q$=����a��f�szJ?좨6<��/�dk��Lj������ҶKZ;�3��d~4&�u��e�^�M}��Ar�ql�y<��ƶ�Z�`2�o�|�%�<Bۺ:}�g�_�1�p��w���k����;OϮ���H���݇�	��9�LLʍ�*�Zhg�I�.<���,�	Q�����_���@�;���^g����ޡT��/т��]�`���QH"�}������mV+��5�"<�)�{��lU�d�v��m��z��P�H�;�]1�T.	x�`9ە7T�ў���@�C�����[���h��I�ה��H m��t���-3Ѡ�_��~tN��r�G+�cp�3dT�'8��Y�������4\�G��eB�)�Z��O��?��D)T��=�q�o���~֥*d6��#�� ��maI�P�����w��T����;b���"��6V/m�H�	l�
EE�	l^�L��l���DM��x���)�N(���W]�a?*`���a�2b�>)�\)����f��F��O_|h�k�������sܒ��Hɣ�+��7��1��w���T�u��������1�pD4,���"���&��5�Ro-С?ԯɼwq�@aR��7���� ��-:W�����[��.|ӢY��?%a�.T�j���2P- �\�ze忼��Ӹ_ԭ9������d��W[�� �G�\�:�~0��q�Z;�b]E*���"g��D����3�bm�^|�
ّb%��'~
�h����Y-�<�~�+$Ut�T�%%�ؿ���T��j�ޯeJH��98�l����T���>C�q̽��)����W,��x/h�Hv�E�	1�(�;:Z2�T46 �w����%/�l����)�W�7�?Q�Q��b?�<gG(5n���UI��ͽ~���Ͻ
����5�1=5f�%�*��_�K
���^�>ova��0\�_WS�*�1�]q?�,F
n�іJ!�}|�
��ˤ�Gb[`p�Èe��݇\#�?^��\�2z�o�mO3��$��lJh�މ���W�;��O�����Gc.x�Q����و��+ɪ�u�j�@��J�y���� �:O8�yҿ�ZK �3Bf���W!�-ea�L]h��5D�m#����
Ń�_��|�r�Yw[���� 9��[tS ^@���)��b����Z�z�=�ß�&N� �6��=ԂҾ��d���J�y4��Bet���;�0Wȱف��_HRM�h�X�%�l�"�rB�/W����@%=�;q�#1���g$�~_���n��ǩ0:d�X�_/��HG�Dy�| �'=l)����#=b#�2��
�|��U�E�v8/��4l�Y����Ѻ)�7�yYe�~���M2x_� 
M�pé���G��_,���^z��c~[�1�`��w�`�����Am��p���R<����gʡ�Td,u��o[�*�,�'J[Mwǯ�E�}5V��/�,����^�_zf�[3MS��Kѵ��;�&��>���fF��ݦͭ�����[�&T���.�GL6��� �4����j&��*LA�Y�:�$��x�T�G��x�S�[�9҄����}��pp��Z!������瀬�8��C����<4�Wqq��Ƞc`�lL`�g��;�gp�9Jv���ai��t�#�;ԀT\��o�r���B�qp��)����ksq$ƃwxB#eS�lW��qv+��W�����D��[�j*V��J ?�p)��ۀ�)�*{��4�^�g>���p�k�j������$;�o���4�g?��S1`��4��Q��#?��A�@��-͞��t��c��LOk:N2���HߐQ�s.�%�w�]����
:Iع:��U�p��c����*��%3k&߱]�f1x�E�<+�.�Gz���6�O�� S����Q�e��@��������΁��[��Kr�tN�;axb����~o�bq$1�R�94�j{ɜQ|},2ۘ����N��{���{��3(�`�͵Xmo\by�����p��2i�3�9d���,ip�na�8^��>���hp�yF��faJ�E��ǯL�-�]�(�I��ތ+`q}R¡��������������ʵ�Vq�ogm{J�>�#a&����lg��o��H��E�y��I����eF=:����2����醃x&2^��*�L�WDq�>z �I�"��j����\j>r���nl;|�9�W�����tc�J"we�6��UzG5K[ķ`b��yTW�5�	f���%W;����N#Ĉm�ٯj�Eӈx�;�A�V�
1�u��W�����Y4�����'�,�!!����a���D#Le�&i��W@"o욗<�6�r�`��*��mg.a_p�!���S�:7�ҙS�]�8GI}��ʁm���F�����؈JdM����7�\D�����^���##��}�`�>��<���G�&�����v����
F�Ss%+C��RW���Zߊ
P��5�f�,B���k;�>:����w�Z��c)�U`�G�	��o�π�W�~Fn��n{��"Q`�PG[2m�AJ++�����ҋ�xXz���T����\�q(� �8�x����Wp��0�-?�;�_�j��ŝ柼 ��(!7��d������y*�?�TA�V7��ik�K�E�+e��#M�
��̕���ǎ�]$w4ҿ��e�hC�M��+�J^T+t�Ĳn�r9ž5JE<,ju��`�t���d�j�L��j{l��v��rq���@/�zД��N�L6�zzF0��1�z�'q�G>ccO���K��x4~���
/�pQ�K�����s�I�?u�ꦑìl��ԟ8Z���4:a���! �͜.k�� @���rE�.��:��;M��D��Y^��5���]@/n5�4vj�5'��6=���b��"�˼�v&>턮��	J��s����;�p,���CuMD������ݙ�~Xk�PK]�v'G��eF9�M2�j��YU�F��F�G9fj&��˄��O�ղZȊ�;�R���d��n�f���924�Π��L�b�n�P����>��93�8|?8G��m��Wr�a�F��o.�c;.�*�NMI43d.���X({#g��&&Eu=U~}C?�|��ܗ��(-B0u&d�O` ��u!�mE������	��h߫<Ә�H:�����کBt[���bu��shd�9z�C��U�o�Ə�����qv*Jh��:hm�E�,�	�C��t�����	�-⋤�Y��o��=n���Z},/�
�I}��C��J�x,��Cp�9�,z�t�,�&�̾bA���G" XF��H</�8{��;���J�d
P7�.���C���6`�3���ˮwy�=�,�9��'��>���|�J��ț��*���.�&q)�a��&�d �q���c8�Ћ�� ���!����7���$�W)$���� �|����h5¡0�~W����A�ND5���^p�z��y1w\q�Ӯ&�5���?�()���J���x4 �&Daď�� G��İ=q�������3��\s�6}ν������%'��wK�&�8xpK3ǧu��O�ѱ�*���L�"�X�[���۬�%t��4N��!�6���V��ټ���A��@?3xF�~@��#<���]�%���b�5};�B}��.=Q��u�=�2�;06P��2OwS{����vc��}�sF�M�Yvc�(���r��`������Z5����Z��T8`n:�A
ݔ����r�r��n5���ja2'E:Ѝi
ѯtS��JT���X�<k����Q+v��OH���rmѡO��MO�:�؋O���g4~�A�"{�V*5ͺ�p4�I� e/	�^�Qc3����@����S,X��L�/^��7�qq��PHS�#zK�eFAKqZ�
�SE� �gj��Kȸ7:�r�i�#�4����Y�ӿ��X�>�U�?d��#h�4�#p��p� �k"iI��iy`�hD){��}���6��ɦ'���[���F�@\��W�'m�ĝ��x#=�:��
��e2�^�h��!��HU0=?K��|�s2hX���5]*>����W2[��v|�h�y�A8n;b�1w��v�k��AiH�<��p��3[W�K��b��w��{�1�tCˋ]YQҪ�0a�꥝�H/�q�Y��a�!���Q���GJ=$��`��x�`O�w�5��@+㾵e23�ks>�uK���Aɮ�Y��s��{��pEq5�����g�*�5�U����eo�tԖ���i�Qo���[�U�,U(�)c�9�H������$Z����{�����ƹC�ZE��xs��0��Yy}����E$���e�,�XYIc��m@; &Q��U��m-q�e�O��4���EH�L�f�N*h=��|���:��7���4ƚ���T���PUL%'��T�LSLY/v����a���^�C�O��+��>�1)le�ۑ�G��˳G�8�<9 �ƀ͜&J�Rӛ�	Z��S�Ix��޹����.�'��y�s2Z?��.w�/sK��_�L����>��ؔ<M��)l�+L����3�ᄜ=�Lp�k��	_��h�0I�&�|��F����f	ɬ��EA��$��鴢R�]gF��������K$����ؑ�H#4"��1��|��Q����v{ L�!�D�Nb	@V�����U�֝ߩR��$�Q���0`HZKuƒ�X��i�v���
u.�\�k����bP�4D�d�f�oR�0��z���0p�m�/���u�dD��Я3��X����m���A�L�6~"�f��d�W�ty�_��(��MgF]N���§���Cr��|���>8���[�l��O�"ollk��R �����F����ũ��
C�/2>:[����r��H��`Y,��8lR�0> �_-��c-O�$@Y6������H��kG�O9���H��A �F{�~�Ithh���#ڗE��c?̿��x���+Yy$�&4�Dڊ�����ؔ��P�?���R9��m�:��g�v*���o��8�=���.�u����&'�`G��@��	w+έ�U0_Bο+(�r�1I�E;�Kz�Z+u�K�0&厏lCK�3!7w�'��C?�|8�lp��D�{��J:�b�W��G���بK>V����*:T�ۑ�v�I��=$��2 N�0l%�\��!b�y������盎��+�b-{�w(�t`ց�J�ʘn_��e7PaӅW:Y`�����gL"IC�u����z[�=��;�=Kf���W����U�IM�,��$�(���\�rY�oӋ�M��P�D[;�8�,m�6�o���Ħ�I&���?
~�u�-a�LF)�>�Қ�ۂ�ɬ���g�8kǮ'l	���e�"_�
��z��X�p-� ����.o`�%>毠`K3���&�3��<�Dy���4��������nvL���vzƂ�(�K�����	Bo�� �sH}����x+���q�k�������9�D(� $O�Rf���3�-�W��;ȼ|Q���Ӧ3��b61��)ߏW!¬���j#6�0X#U��ˠ�NuK�9XQ���ß����������.�*��/R)���i�fI���Jf�޻$�R`���qr�.�Z0�_� �QV�q�0��Z�|�֣1�X�(�u9��,=�wb�c�c�$�\���¤ �Q[~��¿<�p��nSG$i0[�`[gZ�	��ͪ[+�w]�@�wW�����j���cnNJǆ���/�H�R������DS��g�\e���qD��z������?є4g���� �I��4����<��u�I�#��i���eg�A��$�á��aŸ�+dO�*�� �1�76��5��dFP6}5����f�nN|]�A)�¢�P�K��hR_"�
���%����W��2(��H}v�@��nX��VJK�Էk��"{!>�)^B� �X-�D�4�D���=5�M9���#�G��~��)�qJN��Bo+x#��������#��^�ě&�6\U����\�R~Ї�V˅��5X˯5��sK�vGf_~8�m�� 5���-���=�GP�7��L�'�!�	`@��7�pw��,Qm:d���>.!#O�i�G��W[����y��ං�y�%D��hc}�i��|��g�R�vM�B%����U�,�!�ruz�n�E���[��R�;_�AfE&㢌7.1ݩ�"w%��(~�Gmv
��v.�/P��q �ʍZ�p�w�a��k���V\]��1ͩJ����pň�ܪu����1k3�W!�Dmц8<�E��=�o����>�3����5Q�[*��4yM���oԵu��gA󉤣�j�s�"���	�+$������+L�4M�#�s�m�e�\�ώ����#~C���F'>��Z�y�2����$޽�h��q\^�������ܗ�B��J��9���q� {�e�Q��}	.��*L� �S�����9��^���{ ݞ��r6s���㚚)�e�jI \� ��1�������YX�T�&�ʡ�h�{��c��$�Ql��z�(g{-�D�4E�N�ͦ�1�#$���)1��+*��S������ϋ�q�8M�qp��9��d�E�T��aE�o|�X���/Ӂ�縥���K��Z��ѣ]�v�S�$��=)���K��g ù6�l�����6�Kh~�����=mN���}#T��?hL��X��D�V�pFA�;D|�4�TBU �3y~����� 7pE��IZf�_c���f�����Ȍέ�fn����x�� ��g��s���'�]�'�	�>�Vhs*果:�e�����(�p)b�̠*��d��|��6��6�5�xӎX�22�����|�V�J��\���6��*��v0lk��-�s~��j��=Y%X	�EM}����q�������v�ʝLz�y�ٸ.�ϥ��]s�v��z�fU�;As���*���=�����~�������/)��3�hW���1������!�`��)�����ATҩ�1�W2}�S�<
EG7
�.����	��)��Jc�Ng��w�5�(4@<P
ha�Tf����KrI��Q�W-����w[�)ZU/E�+zW���*ўq�v��:�\�[N��|��!6i7�L��I��@k?�(*�?n�q ��jZ	����7A"1Gb�Y�@�
�uj������~������k��%��>f"�W�Oڟ�~�v��[G��#�<ݙ��=�(CN�Gcj�Ɋ�g�L ���G�l ���z���;,fb�\h+��6uJf5&|�t��Y����Jٍ+[���akhk4�i�"��}�ysp!��ӧ�z��$�P��*i���ՌҦ���
��t��a	�o�P�mB��eF�T%��#�9#��w������@;�
�\yh�K.�Č�O�<LX1M�JL(� X��ghR$�-Z +�V�+���1O'���vKZ���!���e�_K��"�5)5���}wdu�*8�c� S�ki���h����n�����<8%;�B���w��F���cd[�M[g��Z79�d�D0��]�]@��.C��b�s���mRD������(��@O������z���4��Ҙܭ�x��_���k��v�P�em�!0�YG��ܣ$��%�{N����DfU
��W9|�S�M�$�֏p2�?7,���`�4��M��{�8<���͙.�4�k�q���(�u�n�ś����qa�z��Q�O=n�@�Z�	�G�ؾA�=����VM�O�{�1,��9#��gb\��Pv,!�8�Z���%7*�M=��^5+���	�Hb���;�¹5�X~5[�+,ZZ��	��C]C�C�11�I��q�r���M�`�)�U|��%G��1y�{�V�ݭbR#no���3�k�yh E�.���`hI��3����dݫjt)-']������n���n�¶s����?0���`R��$����&�G�Gύ��������6�º�=�vC�i���"\�n͹��hR@I�=����j��%(����i()=��}iV�����r˺��{nNx��Ȯ��Z �<�4�Z�� �G�W�ҫ�?p�~U��k�zƝ�P;͔���ܶ* �( �ǥ�:כso���H7&���e-�(�&��'�&�Y��g&(D����������)?�5��xks���H��M���w�TR�z>�CVP�1�w&M�C�K���R�[�SE�PNw؜H]�t߄%iQ��#5���Z1�z&\k�+<M=��j��ĠQ���{�6�Ϻ%L��r-F� ���%8!9��t3�������P' �<���h#�RJ_{�֫�h��L�U���A���)��lD��Zo��o��vT�0-�l�$A��ZK�����!��Z4��v�
Y��לN�n��b�"���Zd�f	j͹.��y�ҥ�abҮ��=��}錺p�� �	�k�\pN������{L��CC�����3��V-q_�7y� ~���=�N���US����7}�h+�1��M;>��,��/�#�� ��qkb��}���P,�q��j�c��*/��kv�\hH��$����3�7D*F���s��ӿ�WU��Ǚ:����Wx�M�ۧ'��4!��c�f$��mGY;6P܅�����V�>�~x�����Mw��3åG���/0�Eo �b6��(j:yp8��2��a��7����Ɂ����W�嫙��#�>�35ڶډS��33�����P�\Nq��o�I�x$yF-� 
$�1Da4��m�$W���^>���x>�o�����b�֎j.sC���`�w��볤5���m~��̼{Mo8�O,7�sZ��	�b�R�$X����h�_Ұ����_�z�ȜGo��깪TUn��G��Ys�1��烂�-�L�rZA����Ar\�@uHD)�bۯ��f���2{d��=4��0���z`���g��ܘu9`��!߯.7@S+Ooz윞�9�iFSt2V�ٽĿ|��}��:��}�nkl� I_�-�<�Ve��̮q� 2�	�R]KA�"f"AQ�E�$�4[�
�F���%2���ϲv{�O���d[�
���V���+�	?S8c��hq��)��DOU)�WJr\Ej(G��� �Bqq�R�QR�ڽ��ǅy;�!m�I����.J�0���o�n�}S�E33��=���r�m�Ѽ�0��EH��ۗ�q=нg�Ɨ�jj��j�t���>��D2�/�3�ۜ���Us�F�/��E�K,M4��Ldka�+�.�/�S5�,����҉���T��ڇy��5ʤ�(���1b���,��}�^8�w�d�*:��?�p挔��|.jlL��Z���Qn�}�'���+��[�Ĭ����x�G<�P�'�aj&1'��L��+b.�|�/Vs�n��E�u��D^��'����&������*�7"b����r�|�[��N(~�"`9�/����ͱ�n�����iO{���ju��[]��v(��Ew���3�e�u�a�]?�+���y5��T�v�ޏuҦ��a ��~���f�>R�0R�>�B8��?:�:��`7�e�H�a(��,�%c�B�i 7��M�yV<w.��ǈl�I���
�,8T.أ.$���v�e[�h�I�֡���c��S�����-����܅n�Tb�bB�m�V��s,y�M���[�r��X����qhِaH/�����L(��T���@��!��2��X^�O�nX��4v�6T��V[��g���
�f:P�jp�Ql���$[j�D�/�/��V��Rw扪����૶>��e�'a�+?�|o��h��8D����=� n,yZ��u<W��bl2��Ʃ�f׵�Z�m��ū��~~!���471h�<	mMćq�20�<�����fE�[ޒ �;�J�տy�1)zᑲ�L�vJ�.����7���$��ڠhħ����s� �r�/�T��3����uÈ�U�X��A����>Wns��˶Π,Fp}�5�l
�Ƣ�8Z�{d����Y����b�&�MX�bf��uJ*���)��&SS�|h�uצ�완�	|���u>|����4q�F���S���b�7�z�
-��d��q�a��5�Q�;�~"=-bA�"f�.�_9��ԗ��������2���\�@:"�Y�-H�ICՅL����,��S�6-��	ld�H�s+=O!h��7����?8-��)�`�S�⻝|��o��k\�[^^j+R�[��)��������]��P��BF��b^��f�w)!rLG�L�
@����&/(�t�-��#�r�}�VQGc��N���K%[�]q+թ"���_��̔9�p�0���ɓ��h������G�2fF��1	�h���^��E�Ky�F�
B`�ł&���.�O�L气~%뷊�,�5/m���sNzľ@�A��ǋX<�>������ߥ��BNMO�eL��Z��۪=�z���wL�b�t��������.}Xe�%.ISR��$[$���Z���v��8g�P<:&���*���"yc��(��I��8����ݛ�Z)K)
�%0Nhh�{�H��B��#��{��8��ԅ����]H^�
c-Y��$�a�v��YD'�gBQ2�����c���"j&v��9䥒G��9��Lʰ��}�(��m񭡷A�􏽾��ǥ�N��~�Rf��.q���^��c��Q/.��o~Vd"�|���ـ�@���Ǿ�K�Ss�ܣ����>%��Uv]�Øri��'��^+�ڿcB D�6�1P������&�tnH%���ɠ[���FU�K�'���@|���5d�/��;�)^_��q��+�p� �0���=�_��O�؆�5}�9Y��n$B�p�6��C��9a7"!��0��+t.���p����"�E���3^ˮ���ˏ[dp�����W�)(E�B��ƈ�-��>��CR,Ѩ&��{UiLD*��s�4r^�D󾎺��%#h���`��������Vص'�/��A��|�5en�:���������Q�b3��Y�vƅM���e�Z.�7��0�97�"iĆ ��$�k�缕��8^�2g�#��/�����ԔG��kA,�(O�Ptd�,�Ο+Y%Zc����sL0Y)H���@֛a��硔�ޙ�l��~WGg���!�S�~c%��F���f:̋��ڱbI�a��w�;��#�����BMg���5��mL������$��7��	�<��v�еeU���	6�lV���йD6�c��#��7̦y����s^��G�a��W_��x���W�Q�3#�m��X�4&��F��S�=W8�C��h}������/t��{��[4����l� ��è���4}����+��-w��H��a�K� ^��!�%��C�q(�/H�q�?��mY>y�U��%]'h�O��!Ț8���u����C�
�,l�纘���U΅�"j���y��p'H����&�OT���q{%�Mz$z������zbV�ba�.a�sphyQ�Vƕ��	���G/1i��O[�1��ErMo��#���':����M�>eˢ&������,:(�՘�����O��e�x�_@���p��|_s#VL�]�!��Z�"6щ=m����h��{�a�S=��*����D6�b#��X�(v���⌓3x��T�������lW����It�]7����d��<HI-�z���pJ��w�񦛀Ģ��V�tg1�}��M&��ފ6��Ԟ�Y�W���];��õ|���P^<ve�%�����?
���' 1.��@��ݭr �ҫ^l�����	5�ێ7�3w3���~|���&�Q��#�,wQCҖ�}�"����Q_c���(�P�i���u.,Y_b	���	�];��ꉐLB���6�������)�z
�����RP�i؇�o9W��������q>�ʪ`A��Ō>�A5�_L��<<�_U��3�f-�Ni��ʽ����/<��۲m�(��w�^f�s���Ov{}��(	b�7�l,�$��6��kV��[\GO�c��$��p��q���`�H� ��#�hM�ֈ�q䕁R�i�����5����Y姛˄ɚ�d�Ǎ^��'�pF��z�YK�73��m�u7hZ�� �1�A3m"�ḵ�����lQv4�x��9X��v4��3�� �*�9��� �1�@/�Q����ԝ��n��N2���!�)5Ǥ�N���a�(.�~X ��EI=�1قݿ�mc|��?zV�pZG�B7�tP���'9�k�Ja�]c��Zb�3�<� ���q�ފ">c�<=?��b�u���"X˧�hM�"�`Ϸ	�:��/T�%%̭v���bpQ벇0��S��X��}��y�y�niH�Y���{a��Y�P�*��%��˟,ǟ~qA0�J�ǘ>��(����R��7���L���)��d���D�|��3�m�&}�A�����3}|�ʺ���T�{�M�<~����E��������N�����叭#�Yj������;�+^~R�8VK�����?���S�bV]'/�HM�XC,<N��"��>/�P]�1�Y�f|�*Tp�Nћe�8�U�Ҷ^��5�(;���� M�g!`�zd�:���jp���?�!CDS�[�↼)�ȑ���MfC�9+��}Z�O���cp���Y� ��G���3:Hl��Z�������$RAcB[s�MU"?��+���bS#�A>�G�km�sZirωzBO�$g.-�����B��fJJI�3!P��1$.U�U�P.'}ց�es���Iǿ
)���,�`�K�s�s�%}wN������~�8{"����˧�g͢��&��|
7����lU��2H�o\�.t�s$wݭ7U�*˨�4�n��׵j
�4�g��pŦ$��"V���d,���M�!t�̯��\ku> ��^u2UB^e�Bc�퓺� �C&g���������Frڎ��|Q�wrN����X�zK����(�׹����bqG��fZ���T���-i�M2w��Ip�z/@�P1��a�LʰԀD�q�
x�L�"tu﫝�p�J�_Ƿ�������5˘܂�c��D�A���������IR���ar,�����>��(ɷﷆ��e���T�њ�=}a���!Ƌ�їs�6O�:��j������a/?W�� �NS��t������.	j���⠏�p�4elZk0�;:u�xj�KaNQ�!6#�v/!���Q����ւ�F����T9�5f���F�獪#���Ø��]��˿W�����-�7Fe��L��w��Eߢ�}��q�2w#�ڈ?��b�y��9Z����a(�U�J���/��{4w���G�᾵K(k�D����#��F�8�`Y�t���2w��b}8��h�2;��|��I}W[��cJ�����V�I�ĵ8ߧ�kZ�MȟМo��ɷ-�M!QmقF�w$5�˫=�ȏ;3��3�kw�'8Ѝ烞wk&KU>ڻ�{!E*��B��r����R�w�$LG>�V��:bhU���.C�vv��/E��A���Le|{vT�s���^���{�CSkַ�-M��ܦp��ʰϓ���|�w�眞Қ��Rrw�\(!�Y	�SN�<�أ;����'ǵH�[�h�P�����c�ۓ��vxB_���Ņ�扖 ��[�:,C�UZ�ƁkV	�gIg��6��ꮐ��G��)c�Ίdm�g.l�Ҫ�]gnA�7n��0��A@�t�U^�>���c��9p��d��BWԎ&��_��v{���Q�	T
�f/t.V��j�F�͌1�/����o���j�;����7� ���.��穸��4U�@%q���`�Z�m�`�XZ�&R�{�I&@�x�;s� ��="�,�;#p�v��s�nu�V	^Sb4�RMdOTCw����R�G�"Y�C$�_�[F1���o6{4�I��y��"���{Æw�/�\��Bq����y�<y�C�#������Y�A��q�}g� F��9X�_"��7�ڞ�K?-��+�Q��X٭T|�Ll�D��q�{=�3�;��#�R� ׶ɩ��y����CsN���'d�z&{3�vĩ<��5ߎN~m�\M�R��k���)'Om��w?��"��$
�r[!���w�ݹ+���Ɋ����q����y��K�*��:0j�T1��!�y#\^�����u{F�S�˚��c�ڣE�����O���CS �?�s�|���V$����H�����7"UC�1Cx^	oX؎f�$m`m�<��h���Y���ށ��I�I��M;��~LƲ(`�r0ځJ.^����s��V'��=���4a/^��Pj��'u��РX_~
�)B.hB��4��lc��B�-�n���'P��: Y8�]���3���ܹ��U��k�r�(h��	�(��Ai3�Z�ԟy �º�]��e��ؼeW���(���g���t$�mv�^�w7�R�^I�������C�un�k�[���HHw�q�#9�;۬x1�N4w��>�)'�T����}Cxb��^fq8d��֡ =A�}kr��^j�8Wib5��y�PA���Pj�.�c���X h�Ub;���E!Jި 6�?��/_@p�y���.BŶ!����"�6U�6�Ԇ|���d�ׂz��Z�����J��p�#�B5��,��=RC��KШ�S����ބ�*	��
�i{>x���Rf<�T���4���+��!c  �i����a7'y�W9�L !7�ix�Υj��8W^;ԐH0l�����q����������:�ی�Zz���^�K�خ��:'떃�bơ���цMv�,9B��.m�2�g�܊��B �+0�����mg�Ӷ���B3K��˱(iDA��� ��	@oE�Xz<�ĞLNd́�s�Vڮ�Gl:��䮓�,�『�ESs����\2��J�.�03p��n��?�cW��A�~�?51�B����:I͏���6���^�W��Q����e4�O+����$\�q(��=+N��R����&0���!�P��Do8;��~���fln�����`˘,�����D��o��<8\�W�����xE����cr�N^_�!��N�����1��8k�+��B�kc����3ي��:Ǧ����wB�$����.B���֌?�S����cֿ�t�	�7����\S)C��!_���l�8���l�26c�zz��t��:���~;�P .)���%j�^��.����>�����ۢ��f:���3CF%�2궐�x�%��(�V��~�FM1EZʞ�dO�Y4�#�/���d&�������{ G����~�-����� ��>g9��.V��'5����"#:���Xޢ��&�mui����]�����A.�R��]M�cR��oΝ�I��M��ϋQ��RQ�=C�իL��^G��u�'&��k+q�㨲Tݣ3�Ӆ<6�l��}VY�X�� f3�}����T\%/gL=��ű}GY�'j�匋��tQ�:l�[���89w%ܩ��i����Q� ����Thu2���N����L�	laZ~��3�S�9ۍ�Y?5A�}�e���G��i�G�G�<�ogt@r�U%@�9�)�r`��VeI��K>f��?^UT����V�ԅ��lv��p�)}n�\��rO����h�~l6��kԖ_TxU��}��?Jrq��M ���uagz���]�ƕ�[���U_@�S��m�xN�$�����V������N�� ހ��f9ݬ�����י��	��֊eX�})����u�o�w9��I��H��C�r��g�j���� <6w�S�ѩ#ĺټ�M�{i��m90L��G>Y�
�G\++������a�3�](�].�"���#�F�t}U뫝E�iƉ�U1�b����O��o�M5c3
����$�g�?F�L�K��?jF�׫��.�t����� Y�,������=���g�}ʝil�Xj�\a�A*X�K��d��=yJTJB2��@,�ccnh
���e�ܨ��7��E�W���ޫ>jSLX�Zj�|b3�_����Y�C�D�(N���+�ϸb/�-�}���&�P�>���=)�>�t��n���ױ%��,f�!��n�''�2��đ�ìR�Kf���
/��[B�� �E�W�	c�?ko`?�0��K�e���b#gs46�~Չ�3����R����EF�"ײ9I�Q�/�:�XS�e��2�X/GHc��QK�X�{�iІQ$�����X*�8�5?�}����k%�.�V��O��[����B-Ps��Iɋ��AM��"q:ȍ�p=&f(���V3x�ѵ�l���-$VhR�4_(�"���Ƃ���!o�A�p�j=���@J%f�عx7�G.,��j�7&8��d�I���:����
<x��21�+i�r�%VD���s���g?���	�#��� Z}	��[�9�ar�㷥se�����Lq#��I�}�k�n���f��:�	�9���P�����o2�}�k�;�=�DQ���)���� t���MZ�#����5Жr*�n�d&�i{���6j������/ kj��	�,�����WǦ-<���|[Bʀu��s��S�7�پTR�ky߆Y�)�p�m7���ӖHw�9��>~4T9��XO���o,���y�lmqG�eHGCtG�)�V'ۿ��Ö����41��S��nFޅ���!���@m��	�b��R����>���j
�Ǐ�:LPr
���	ԗ�#�7�ro���BB����)3�i]���bAZ��*�܎V%�7�7�l+�\��u6��z%y�
=�.��Xy;���BfI-���5�Ӳ�W�B�:�s��/J�}k}9�C.z��`To�P 	�G�0�S�Br���'i�7��Op�!�7z��>i��M<�a\�e�����gCꈉo~��Q��1��I!���y�#��U�kkg�7%�U��I_3٫�H�ݏfV}u���8�TNJQ�����0>;�S4h�aLs-���#Ugj�_߯B��U��.�D/���@N����t	�ZXgt���4��*,��2���<O�����
����`���2f|{�>���h�'�{qH��)�Ӡ�R� ����3��ͻ�*c���D�X��ٝ�)�����ǥ�fa���P;=�f��-�A؉k|�&�b���Ƌ9�2%p%��{
7��+�9�t7Xa�x�$]Q�}Rm ��(��k�s�pJ��Q�{su���r�����ch�Q�{�W!8ѳ.����2��I���?����������� =�E�]�5�T�/s�	<�%Y�a�*�К��ũ �-�yAh/Aa�0	7�0�n�2_*������7��cG�"4�')X��b�����y�OBl�*U��]������{~.ﻷ.�TX���;��^-A��dc
8H���"G�3U���Hg2���]%��ßu HN~�ș3��}m�����,/�%��Y�w�»�V�i�9�M�xs�l¶i��M�E�_[n�s�$sӵɄxˢ7�Ї��Ƿxq$j
%-~�G�d�2�W9�fA���]u����������<�֨EtAMl"�;�s�u��L��z��:����Sq���T�RFbs�}�T�$�l�_=A@�N�x�٪ΝM:OR�J�}��"f��܈��L�jG�M���^}^ʹv�c�e��Wz��LE�e�u��9J�qK��-���ko7�Fl��ۻ�)7��F8�R�.�=s0=��x�W+v�}�ê�J�9&&�~��7eVĒ���2��Z�X qzq����Z�ڛ�N,�������MgyAhr.�H��.�9v;�l����r6�(��6.V��'���L b[��Ur�lȅT�������A0u%�&`n"�4⟌-;)�%J��.�/k��-Y�,]
l󍋀 �m��^�Cp:7�Vf��B��@Y�PU���0�X7��prҫ�����;�y�"wy�7�⚻��::���E��Dm��d�(Q���y�%�$���8|������:%�HGL]g�r��G,=o��"]�M
	N݋bW�ij`����MZ���P��ڼ��7��q��N�Ú'�;@}!E������T�WM�-���D"�����hn6_X��T��Dr�~�P�?W��%��K/%~��/��!�߹�v�'�u�Xf�$�� �����&*g�m�/Ip���c�����Ǥ�o�.*�/#����RP�_�.�Ԇ�>)�~�����j�_(�.9:�9���[)�*e|�q0� ��]�Cb�����7�U�`�n�2:��D��ja�s��Ȉ��)�v�	y���6�������,[�[=���ʦD�:$��pj����u�sg�?�p������?:\W2]�Ԃ8��+��*1���2Ëkg�]�h6���x��r:�B������6>Z߉�EO�V-ȃ"Q�������rGS��Y�k2M�.:]����R�>h��I"�uҋX>=P~�Uzu �>:��S��r�l����8]&�N�	���4�! �8ԩ(�F禚"!k�耎�	&t��ƥ�1�u��W�Io�v�J&�jb�d����x�����|2V�E�uu�3����9(�@�O�L����z��䊳�%)�� ���rH���7��b���-h�l��4X�2GP]���@PCޣ��[E�K�,���#������h�,p�~��f����ކ*�c�Zځ�t�.b�B0�	w8�F��@�R�I5���J�"c=���l�0W��~��҈9��&���=g�QT�*9u����LCz��}�ChtF�׉��VY�t�h��lkQ�0��~ѥ�Y���+2�WW� 0�+$C8��$5E]���܁�z��,���8�gn���+F4HppS�ж�m��}�r|�'���+ն3f������
=Z�]/y��yL���<�~y:Ǐ�q	�Q�b*�"S�	�U\a������[u=\#U;bH�͜�zt�܋�TTF%+w1��m��R�[e��VsB�!�%�������|��L]$�z)M<�7�Im�k�#z)(�.��V��ofH�^��c[ƪ(g�=?�<�8n�9IZ���#��ӆf�s�׵��ܗ�zi��6O�_WݤVm|d����ʝ�=���x��%���[hͧ�87��1�'����������~��f���nKVa�[�ˆ�.r��ze�xX��{�ӽ���9ȧ��>q�BMG�H��v��z��F�z��P���uS�+}<v7��mHQ�f��pF��[��h'\lJ�dx�Z��Ƀ7�~�X���"+�� �#�j�_�����5�6�A����Q"��(be/����u�[�	����S`NU��s������Μ?S�������Nv���oU副C��d��VK[ƣ9��O�e*�4w7�`�Gk߳d���éU^�ۂ(A@HD�U���>[v�~D�]9z�Ҫ���;{a��0�1����c׬[�����LI��V �q��"�Z�5�髿��]����#p�mM����ä5�8�?�!�b�O��;���Ei#lj���ӝ5{UV�A&�
4,^lz�qQ�z���k�?��g+1�R�q(���l�h����+��;��&)�{efz�px'�Tu� #W�6�2
Ԧ��o)��T�;D�S��˔(;O�1̓=�ɍ�q4�븮���Ae[#j�>�f�ϖ�e*56�k �Մ��T�x>�K")�a��7��14�_R����ͦ�I׸F ��J� ��<��[-y�N���$��U��H�������������`���n"	GGzV�N�(CR������u�`�pW3�̤ɰ��JJO��q�Ł�������^Ⱦ����u:�ö'�u�y�-.*�~�����U�WD��Õ�⦅I��5�5���4�!⩖]_�{� :���hd�[v%lm���GNi_v��� ]u��$���ۋgB��+��~�a�[�.���B�D�+qE��[>/��č U���M�ƨ������o�N��:�����A��¾���5��v=�`TN��!Ҝԯ���0bs�,�^$	�?�>�	�GY��mYa�bo�<b���ő;���9�;��۲�߯��K�35J�M;�4d�yٚ�?�T���ȄҺ���>Ns�f�!C��G�l�O��,��� �'����ƣ:�pP�u�+����{�	����ゴ������h�Χׯ��$�`��I�����H�O��~־�����^��)Xn�ߘL���D�l���Ǘy1�EО&�e��jQmw���(�0e�~�U!��2��HcE&�c��z�Qm��[G�ډ�33�w�}�Fޙ
ޭz�pp� �ゎ��Yy�]3 �=���hB~�7�K!'WX������1���� ��w@���7�D��B�K������K�O�yL�P�S�*7��Щ�[�]ófw��#���0��F�� �Zо�=�Ӆʅo�R8�&���9L�����$;;#\�L�12c2�W����@\q�;'�ǪX^T&M���p�}� �ȀD����uB��#�3T1S�����f�p �����H������Є�Q�o搾~ݲO�늠����I��L��x����IC�3��_��
�����wYsf�����#���=���;d^�z�;���	*	a5MZ�r��������,�k�g��e49J������+�_��ӀԆ��jZ�p�9
+X�5
�d��3Ts�Z�TM+I�ߟ	�����;�6-'�n]7_�fp@�6�9��O��Ñ��`6$� �½��R���[����Y���8c_��)�J%Ŝ="۩h�u�����GcD���C�ct�99��e#
ӏ1 8�H�XV>��#��������?Ш�V�T���������3���y���<��0?\���qf}�9�t:���g0_/X��V�c�u��_�j�T"S1N'���W{��h\i�FȤ�.$5_y>o�vՏ�<��p�o�0����od�>����a?k*�Qi��:~�qD
���R-�m˙��)T�Lό���>��V�r�4�`�����7REԫc"Ȧ�ā�y�E	fOz���ݤ�l:�����������}�|�u�c#(��+�Ŭ9��H>����ik��!�綴�~wڜ.݁eRQu��V�x���[�A]��s^�D���[MY0����\���5�����`x*m�n���M�\}5Y��.]_g*�u�8םd.� �a@�-'Y<@�D����AN�ڄ�r�ٗ{[�J����^�H�`���_���W;�E|	f�1�;��E�Qiógw>�Qa\�=R�o4��`�~b�s�O�N}r:8ct�����O��!�L�+22?�E����_�,���Z��CS�쯡��,g���o(En"_0T+b+H�g���j� ���fDލ�N�1�V���/����ۡ#�pqw�3SW*�\w��L:�@3��� ���d�[�������ٺ��=��l�%�s�_1Fr$�Ԕ|��j�υ�E�D�C���f��G򢞇Y���=��T����fs���$Ά3Z=B�7}`7���]�n��.��(%'�篜�Q�h\��7���]e��Ja�]�FY�S��,��W�i)��L���t)'r�K��@��b-���Q���;�P�N�ޤ�\<���~b����%ū�~>��e)�~�r�9C���xƙKk���r9���	ѳ��Ƽ,U9~�gJ߉�1+$���3r�{۽=%b{=`ƅNI�s=���J�]I�P�	ڟ'O����[Nnn'�'���	����Н���ƍiɝ�_�-O:�@;-���?	s�霾鳗����_�`�>o�	=QI]�h�U-�I����҂���40��Ȅ�|{v�kat�!j{WA�J]�?RE5:���7���P�
�*�Hk.(Z[1���>�1%n�@k�2A^^����'��s� ��+ff`�й2{�Y��g��HW���׊d�n0#l�d���h`�O�]�݅�s9>��`� �8�<�v1Tht���L@`ު�vSDpi�<Q�o�?9_=SCGS�ym�A���s��$��@�a��ב�O�-��5�q+�H���4��՗�!:D�PK�� �n��Z�������&R	x��O�)��T_E(m.(F�	���
3"�jh�3�aB�Y��]��>�F#lC(�Fl��4I��,H],ث�$��	S�pz��Z�
�
�_R<�ݞ�5����5r#y&;���UL����rM;����M����(+���%ק�G��?u�(G9<�a�i3��
1�NH����ī4Po�w��w�G���̙�擯]t�`8�>��,^��-#���5v�^�J�lI��p1�j�ɵ�
?�gi<���o��9�i'p��g�J��Kn���|�k��V.��~����|v����\�3t�Rǅ���j"�Z���S��2]��js���$��l	���ҿ|�F�A�x�-#�ׁcȻ,⍚��d��!De�����f�^�P��qSk�'X�=��0�,9��j��K=	�
�:i5�{�M���
���)�������Y��A��wv-��)�Ea���B9�Os4EG)��q����Hû#|��o�F��u�O �� u�}��Y���y&'C�������#9���.��+Jg�w�Qⓕ�M��	����:N_��,�I%�m·��}.^���1�?
ohm���ՠ�S�"�~ջ�ԅһ$�'���B�4-�'UƑ#�ճe��d����m�k��Y�ҵ9�
�l;���g��z���B�s!�vjUǾ=��}��-B󐪧���RU�a~��e���"*Rۨ��6�~���"�h�8	hC������3�nm���_��G�F�A����>�i�v?/����׶`�Q��!W]:��������9��a8�u�L�(?����v���87��в0L1�B��ZxM�0w'M����U�%��M�rT1�[8=[�8�wl2'�k���f�4S�m��cq�ff��Uj�����I�g�O�V� �D�/Yg/o���L� }���n66�-1_xE~}�bJp�H�Ef��#�����u��"!z
���'�x��۟��i�_n|���5k���j��.�ܒ����:?�H�"
Y�xcO��xȂ�(�Mk�(����KT��)���}�kf�K�gU܋����	�Q�{N���x�<i4PtMr�4���C~�ιH���H0`>�{!�_�KY�#̀l[�{� G�5���J����7U�H��-Wo�
���݋G���|���x+ZiY����-!]Ji�$�A��6G�3�8�oB�0K#>i��~;�g���՝X�}W��?S��vӕ�c^�R0��ɕqd�N���4�Ab��UE����|��Q&� �=�E�P�6-2�!����xڱDI �@9�v�
�D��}�c���Ӂ+ �ވ�B+��,��s��qB��U��l��4Ւ��M�/G�G���ͤ�H��6�V&�
�e�����y�!���F�?	Q�ixП�{G�`H�ʗ?qD'��!�
K��%G&���3�V�r��&C�:��ѡ̔xi�_�FJyh1c�9�|����WR��{]Ph��[��1�O�f�)�8��kG�Fa�#�_��1�	� ['��
�TrSO������hR8�4Va�_��7˩�L$LQO3�ŃZ]թ��\�A�,�(��m�5���\�bA�ptI:��^a�y����ZL>"�IσT��6j:��|��掔��i��?�A4�Òۦ��[���u�����,2<�_t4����axp��{<!��6����{��;����q&���L�'�����?O�`T��ͦ�2��9I5V��MBm5X��DْQDgce�:6��H(Bs����x��ʼ��*�sF�O�.������#����a�<�3�eCǠf�}�]a}����r�>�sF��h`�g���ə\a��P:8�����',�z9�)��.)K��ᚺTv[x�Ed!����o�������ME�6HԪ�^�߈�&G&��.4�y^m��`�ب��K���m���#��A�a���=)�R������zd����ёPV�������SCNr��k _�%�cb�eU�H�kQ�*�LI�*����>�@�ƒ���T�BJ_­΀If�����#����7z*M&e[�!�F��=O#*j���2�,�K����[��.-��E��V����ק��CZV�;�+���"�1�]6//J�ߘ�:l�ƭu*Qh�aN/�f���è����}���A+ҳ�|�Ω�vd��!kNtY��.ׇ��Ɍ��t��p����CMf�Þ�$�h�
>�s�/L�y4�
ǎG�}~ t9�nf�ig�lz|w�Ix!�	�LJ~�T�1R��V���B��~-ܔ$��8��'۹�
�p+�z��B�;#,�&�{9��EG�[w�o���$�Q*�$7�pWj�?qt|1��W��-\2����yX� :��@K�j5��bڒ�kݟ�t�A+}99.��64�KH�vC'����c�p�s���u�#J���#�`]��n�z�HSUo�S�Sh�Բ@�>V�?$<�|E�1�԰�ؤ}��#'�ڔ.j�����ή'F$�b��]:�#}�]W_X��s�t��~���;�bA�XU����vj�v�X	�t@���,����xj��	ˉ�ϫec�o�v�Oִ'�Y��:��02�(m~�04,2�����$�R��,��p:��*�w��{_��"h���������)��f�f��"��I�GiI�;V��ݓ$(4{H%^�ex����`)����������*e��'y�w�h�8���[~��ğ5�a����0�����ľ���M�c� 3���X�ueO��>��M_%M4��bh�ٵYA��cH��2��"�\˯>oW�F�����ϹB�"�1��|5�.�nԓE�~	�ld�N'��]�֯;�C��RD�ӏ���!���}�{{�v �ĺ��	ҡ
Vz�L��Fچ-�.��7��\�Q�]�;�"��ʉ�����-��k��@4�%��3�>%�[�W��F��;T����ِf���b��TN��W�g�ר'�G�ii��i4�:����e�G�ypYe:�?�,��J���y+L������������ŋD�������Y�p��GO�,�́�Q6_݌�}W�S*^{)����j���b��xcߡC�>=�������V����4�r��:E4
�x�M�[�	kt�GRt^�M��f����E�T��6Bb,�ж��.�Yu.���J(����8���B�w��Y����1��j&��~%ߎcٓ���<��ҹ�����i�S�k�@���.����D�Y�Q,����8��@��Iu�P+l�@~D�`>֨�yx\_�иH��#.[��d�Jr&u<�[�a�x�-�?��j�^)^�9D6��d����օ��>#����+Fl�h���_��,<�* ;9F�b��P;@iL��N5�f�VL����i_���=�(;�>�@��h�%r�z��-�w�m^ւ�I�,�M���2�m������kQ�)�i�K�@S���}��#.��]�j�d�h^�X�R�5c���~��eM��#v-� R� ,5^�����h�d�=�Rvapx���j� 	uF+�����������*'&6I�������֧�'`j:=Ɠq�j����lgj41���B�6U���0��A����i��ZbL�mVӫ��9���z����"�	զբY� �#���ʲY��B{���p�=P��_�gO�r9 �b7n�'�Q"�_P��Hed�����3J.�͇�H��x�t�����'0�����0����"�Fqw������qÉX3 ����?;Z�/�}h��eE(my���D�	�&���e�y�nk^g��2��
Z��4���&�6���F��gXh�1	���)��{�o�d�F#Y��bxrK��d`CPP�YoB�:y��oc9��b\=�^����%�v��	5C�D� �ǂ�*'�d���>�D�_�-�����Da'o�Ep��XrH�,J�w���8JM����E��:�O�:�<좧�):B�Sr@L�ݧI$j���䵲Ɇ@�Z`t��$�߸{�ċ	�e}��чq�x��jM��x��,<����D|��b��v���a�?�	�+2�ⴠ��\^1��j�t��}�5}!Ik�ђB���a�WH9w�T<%e��{8|�Op��kY���9��*�9�^��[�<���h��9��%�+������l7,�$����Q�U.��R��S}j�����5�\�jY(��w'<�D���Ӂ����&GL��~
���l�Q�I|q��Nэӗ�m������o��N8����r���j��s6ɚ�N"�{��j/��K|��(�rݞ��I,!z���ݜ*)���}d�����Cs�&N�Z���^
D���Y����AvAB�ߡ�����	��������h`{0F��$_U6���h�qx�j��BǠ������ݓJY'Sζ{��\H��[c�3c�[>/��^�Q�s`�HYF��A��l�(��S⊨c��	��2$4#l���X��Ʊ�)�0�\�c�O�Ѭ𖉀����*��=�}Ԏ��7^��=��`�ŔQx�̂-��e�	��!2aQ)�=j."�����zw�6��N2�x�i�7�����f*��3P/DR{�N���4N�J�()!d�E����F���'g?��݇��$��W���6ucX2&*0��XVf!���yY�je����?���������F�YHs��y��f
f������Kf�Z��P��R�q��h��>��D���{�q0^�����,*�lr��PA*߄
��	���Ņ1���Ύ�q>��J|�e�͉�VG�3������:��O��#���4G�G��êL��������WΉ�()S��D[���z���43�!�6`=y����#j�~&Q]�&���.0c�h�N��1����l9�/>�n�7H =�2���rة	c[��ó�I�w_�C���A �GQG�5��U�\G��s�1v��������2t���f�Ak0t4X�m�^���O�~����
����J�������֯R�*�ՆiQD}�#H'˅���V�O5V�`�p�TD��gp�(���@�|o��t�O8���^w�*����t�v�y�gi�W��U�e�yC@��N�gb-���U4E���I�Z9K[_������g�j���e���\�P�FU�A�ɭ�.-~{��ZO�o��g��Q"0�p��x�M��W�ԝo��700�1���<p��L��8��ݳTâ*B�	_������&3?J����'��x�`���<z����W	�G����u`���]���.i���p�wUՆ�&1���� ��g��@W���u��)��.�>a��E�������̣:g��[��>d���m��׫�<��u�4k��H�7|��e	�@�fj��؈4<-�Lͅ��і �L ��=���P�M�.�]������_���Թ#��}9��}��t��}��������B1p�*7���v>1U��.�BKX<�}!BW��C�S�ږ:B�[���i��9?t;�K�xMF{�y�`�-r�0}m^Ր�}z��j����@%,�u���L=�����OZc]�!3���D��-Hy������f��S���p�;�\/����m���Db8P}֯5Ex�N"ԍ��h�l�}Wp�W��#��|B��� ���yh�����B���5������Y�찂�� u/�a�k��s�#v��|;���=��4�w"�I4^�Q`qq��Q6Q�+
�%��qX,K�(m�|�O��ÕV�m2;l�0nXȘ�vG���X�&����2r���4�E��P� O��OP��$m��� p��`�G���z����U1�
��*��5�|�V�O7lS����$��N�ۻ�ء+p���L�T�4�6��z�d^t9��׸>u���ު�|�ߦ�H�[Y�(˓iJ� ��uX�ޢ��L�?�U���mڛ�g�S��1���zO�\��+�|������MW�8�Д���l�eG��|]��n �ED�A�%z�s.!��N������.h �j:2$6�k���#�Xx�'����C��%�i^���~�+_{97@LA(F���[k���{o�o�_��_��)iI���(��B�d�%��Eg�
sscW�FQM��w�Xf�*���i�r8�1˭s��b7L�[G7/����Ƃ�@��&�ͰfK*�0Jf܁̱!;�Q�\���-k<2 �TF�Iܸ�s��-��V�������?_����<����Cn�{���H3v�U��>j��Z9P�B��/&�A	�
Itp��S�=���-�CĢ�|_Rx׳y��ϩBC�^�f7K�׿�;�OQ�[r&�I�f�-�o���dAG�zu��|89cE��v��V������t-"_�~0��.`�8^W�߂�V	ɓ*���qk��s9�� ��В�00��R��=�|���8bϊ@�k��B�=�Xᦋ�P��Fŧ�ʙ�?d���f4�*$���~����{ .F�?��Q<�&���M���A�;��~�;���g��-w&�p
7�ݛ��o��]96daz���y�}}|(k,҂6J�G�GN���(��_v\�����B"u�Ef�M�,��# ��eE�[�(�u���VAoH �P��D��3+J�[��>�?�u0њ8�M��FuW�X�8���/}�(����������URDO�o��^��e��/S�)��"+�61�irұ���a�i4n���%�h�����E,��/_�|Xm垛㖵>�T]A��H�!��'��Y��z���}G���慿Ht�{T7W�^=�]{�����Ni�Է��~f}:R,�0{�"������
��
I����"����&�5���s	�������b�"�x����&��o&a���\�,01�A��j
��v��6@��ᐲ���j�����ƿ�v��@S�&}���l42X2c4��cYK���d�Q�����&��/���u��D���Ԝ3F�RXiS�S��c�_�K�|�X(�n�c�>W�Z/�k�*�֍���f`���-3nC�?^d
dW_*��$��̱T����Np���o$B��3�C��B��7����
�<s�|�қ�A�>��Z�#� ��Ը���B�b���ve�Q�x4���j��,ě�L�ˣ�{�����Zu�宕C�L���R�����v���ʛLm۰�:?�n1�E�(��K�����9V��P�K��݀p��C4_Ҹf�OBT�F-��k�����;|7w�*���\@j���Y��jZ�BJ/#-^�4�ݘ�G:G�Џ\�Hɠ����U];��{#�Ϲ�a��כ�W��*����(�hd����A�������	���=��l,�e�kz�+�)q,��
���2�J�R!p'D=���EF��J	��5�R&���/9p��i���(y�4��p��F�+��L@�ey�KC�^%��Of"�K��p_����� P-J�M�f�S�w��<� �thY���D���.�7�B	�A�wV���� =�
9a~��[B-��h�7
����h� �k��	��>�S@0��i�~������q>�>Kh�+M �1���̜�c�,�m�&u/�:�[�K�����6H5�P%�yBj�vKľv�P{dwc��ڬ��� �ߓ�?"R�n1]=�[�Z�Fv��ş����-���F�����V������)DQ� �b���pM��Nv��9�;}'�3$s���t�S�*c-*0H���Ip�;:^Ct��n�*~r�ՅTN�\��3�0�,������w{�owZG�R:��{t���M�z��o�+�_��K�mTB)�W+��SPN��OX0Ԓvߊ��I��CI�*��~ځ�ܐ�"��B��~���T�o����]u�~a ���!_	i����{�I%]��=h7]U�$���T��'�x�[ܞ�r�*XS��.�9�����^wETZ���Fc����ɉ�>���Y�iА�fdP���U��GBlZ����y�^Z2ړ	�5r[(F|Q<�gMns�a7��̥"�ϒ�V�k�D]�s��t��y�����c8�sc�Y��w��0�b�3/
�J}h��_��#<b��;��^�e�f��/���
6P�H�L��#�M����ԬT�~!]'JT���o|3"��6z)à�	Yy�=Ɋ=�x��T\�m������c-�ߨ�}��萃μ/��i�����	YS��]s}���M�j��=q�����f.�lse_�q�VTa��C�'Q���Zj4�qYz�@m
�&�����{+���s�@ns�'R
5�ͫCЎ4'���[�Et���+���҇\Yv����<��K�J��XԀM�i�3kI�a�b(�`ġ���R�b^ж����ҍ*�;Y�Gn�Fi��iC�V�����\�ٴ�Q����e�z��c�K�RYW����&���8"��R���b� �z���"`lM48�I@'L�h��^
/�f��}�M�X�h&��$4��q���d�lqm]aXٍ���fY��I�����F˲]��`-��Q��@�fy�����~��[�u�?�%����G0mnKOw��4�:��}~�[q�%	^�`@��yJk�����n$�y�e��E��)_x�}|~�_�ޅٝkr¹��%1�f�J�Q��ǌ>�}Ū�Z YFdk��H<��n��f�$c{�N�RC�b�7�j-��bRj�������}k��V�j���8Jڈ.���e���+���X���>��x��(/�j)��t�$p5)t1�O�X�;���֘<j��Ў�qU%�!�0�Rl�f����۹;��c�?�G&���R��<)7��8J.�]W�J���ĳ�!��`��}�ǦV��T%~f��$�5��!͑��W|-��ri�8��"�?��T�(�Z %�X(a��#-b�G���.k����(��jO��D�����nخQ`TFW�"���S0\D��7D�<:N˄�	j�&�)����>
��%��Fgf�#ĝn/�G�!�b��J�ܘS�k���:C�w~�2��x�>���\|4
R�x��̾N;�Be�T�ƛ!G*�������
]b��5��8Bqc�;���z^Z���I0�ʬ��Dx��Z�{P0)�'��Jk��z�#�B$u�
��9�o'�a9�;�\���`����=5Y�9�7ڤ�Ghg'O��%��mW���n��5`���0͇N��ԯ/X�[�|Nj��H�@w��<�
ǂ`9f��p�p1:e�\,�� ��9ͪ�~�g��tj5l@�&�ض��K[�����6��B�eq>R�]H�/�|��Rk����V�:I�2���$F$�\�i�I���E�"�Wco+6ެ���|R�޳t�
��|�{��Ԥk`n7�L����|`�b�[��?X����j����˪�$V�;��>�H��e�&d���$��4т�;g�!S.���#��);XIGF�k��"�Ŗ��;Y���e1���'�^��2v��!>��!�``
�[^t�u*����s� n��Q_�?MMF��T07��G,�<�!1o�
�sEГE�9��q�2^?�bW��u�A0=Vw�yy��o!ڍ�;��4��q`ٞ<lVZ�Oi��ps>�C�W��f\v�d����H}r!
xD!Nϩ9aH��	.�ں(��D@���~v���%���{�#L��Vy��n�t�6���Tj�iwj��Om��4��nBY��do>��>��Ӕ,i��%��"?��zCG,?�p�@#���w+���r�J����閟��;�A$6�^�x�!96񩇻����41Տ�|]�_&��%�4ϔ�Ԋ\⎐� �P�{��w�Iy�I�|7hT��3Hl��	�vŸs�� ����I��梂�y���~�Ư��l�K��8B�]��7Vz#c�ʔB�LJ� �0����E�qS��[�8��~�t7	��	�P�ܷ�n	�^�ے��.k�X�j�I��ԓ���N��q����6�b�/� @`A#_�Y�ס�;���K�+��1��h�{ ���z%�Xyv�ܳ�J1�ڣowFvK�
u9�rK��%X��ۼчP&r�%��z"�r}U�K� m��l�a�(Xtv}��ʨ�W^5�]m�i���h�6b[$U�r���Y&�4�y�c����˼x��qi��9&l�eb��Z4 BW�Pb~'H+\�U����/<���1y~ǈ�C6�=�=��ޮ$zH��h�4�����a�2�~��Rw��I4)����M��%�N+��Jɀ+�k��ɇ0ZG�'��f'�%=�W)uӸ�M�
��BW��5l-FK������|��S�Đ�#P�m���G���닗Ѷ��*�b���KH)��-�F��w�)l�q���W!�E�����G�r�Ȧ�⽉�zr���춒�M~�������#�����/Cs��+���@OB>�r���z���l� b=q��yњ�8M���6��1���4�[�/Og��qtK�mD��ON�>:�(��c������+hW�Ip�����A���,ϖiU��믡{mix�Wߟ��.�m7���3�7���[�%[Tr���k�mD_xj���c�)A&!�%��ʄ(J$�K%��ֺ�8�vI�a��\�����A��$�c�(Sh�l��I�Ү��0��}�$U�(����Wn�Gj��(ؓA�X���q�������y�͐����"q���rU�zk2��b:-^�@����#�epui�IC�Hϧ���*}�Z��尌U�����<R��@4���ִ�rkK���.��?�3��Nz��Jۥ�=����}3o76"r�˹�m��dC��tߪ� P���`X�L6�>f+U��(��ʦ�%h��g4A�p��<g�:����$�ow:�n��LC�v� �����:z�69gQ.Q��45�
1m�BG��-n�$Ҫ]�b���G���Q�_2�����ȂRܳ:Ő|��y����daOp�^#�%���t�����H<�ˢ�]�х����*�
��l����1�PVUu1�+�لͬ�}�E��R���ȉ]%	���d�	��;���IB����t�<_�Ԧ' ��H�����:�Q#7����Jܦ��ճv��|?w����G�� ����[��~��,9.�gX�)��:�(����ku��Ȏ��	����E󳷥���|i/�R}�;Ue��F�$zl(�P���;WR�? ��L���p�� M%n={��c�	a�����mfÞWiV>s�}�ų��f���bz-��)'v<�sE�O��Ii>㸗��q�@�-��`H9�AN��<�=�pGh1'��*�te�������8�d��%E�NSFYД��T��� ���f���l-be�$&��pj�u�b�C��)t�,��R<)�7h�j�\�%驂de����ɖYǿ��� �t�Z�Bxٽ�<����${�&6�W�P}UF7�iٌ/�U�Z%�����m����ﮨ}�Ć=e��m"��l�3��Ά]~u�������ڏJa���Ԗl���J�5����y͞;����@�}����Tn��dxe�Z]�}�͵��m��]	�^NR�2��&~�ə�u������ֽ{�*���8��s3j��b�Q��D�gS�;2
���0���~ڰ�K߇��lӭX�6;V�6�g_A�e�N+:"T�x	���C*[3���J2�`N���,�y����~!ϧ�S����9}|��|4Z~伐9kELyxg�&l�@9Êܭ�Z���I�\��/��fGꚭ�\A�k]���U|wN���dnbBM<��<���7�T��j�^M�e���O�y�h��V����m�H�ORj��-��a�C�ؽDa�;Ԋ�/O[RA-��C��-��E9�
���S"t��21��݉�߷F#t��6Ȣ2�����A�*JCV�)����/u>I���.�m�8�١".�㡥$k�� ׾�/�d;�*��-\:���!J.��e�ڸ.L��
[�l�	]xf:y�&ɐ��u�f}�vsR��7��g6���SA�����0�	yP�6HA�īlo)�K8�C(��K���eaa�&Zs_�Y���0��ȇb0�v7�JIZ	�(-��S������7� ���l� LR:\}��7�S}d�x�K���V��A�.�޿��k��mE<H�q]��3os\"XX`O��u��*z�y�b�]��Y�eXy'֎�h�)E���\�4������U%p�JɅ.�"nG��z)��ɶiD�A���!��d�b��
�_H�sy���
jE����y�ŽbAY�!"�qԺVV����H3LG���-��v7'
1TR��7�C�䪃쩹����!�7t���=����M�;��}s~!<����(X��zv���%���� �N��Vu%���s�'Ha�b�(u��;צA�7@���1�0j ���h��^	6C��j�����w�ߔ�#�#hV뤚��l`����d�E�;_��V�;���0sv�bUľ��+�1|>���ukfA���X��LM"���XZ��!�Ad%VBW#G+��ğ^
tM�J��&��ɟ{yNi��	ן#����`�T��U���O 
��{��h.q�"�%:�zxe^�_�FԲ�9��^2Q�˙%9����}�pO}��6����Z���]�"}��X|"��4x�ړ@@w��W9{FZw��AΉ��f,��\$L�R9����b�Fio  �Ӻwp޴����:P�f�vaU��oP>+�%��F�jG�1�,�p���@�@#���0�Eٱ-�������^W�(��fO�g#~���~�x�2/3��ٲ�O'{� �&�?G�0������g7��?��dP"\vҲ�9������>D�B�E�-zg9�ݰ˺d��?)!Uу�b��E_!"��W� ��%��O {�L�Xx��b_�s}�֕��#0�,��{!$������.�_8���'!�ʣ��V�Z�,�T"�[�q	�$kdH�5~;��8��
������a)$3��qF�,R+�Ǎv7�9����s�o4�52�0�v,Ｚ�UB��OTm�Kؙzy����5��{I���; ������/ޢU��o����J��U�g�;��w+��$)�*e bz�TG�������ױ�(1��?��_"zR:�m��	n���6�C칝�F���,�����c؄9�?����~'�L]k�����T�N�����̓Cd^b�rJ���p�:��2���R�|�G$mΗ�DB�&�G����ߵ�S��0v�Wfg2�)��uQon�<��|.�C�R ��؃D#�����bnSѻw�t�u:B���r��<�"frf~�%�1��������*),C�@�$H��/c�5m�_�#z��8�	�*����*(:|�¨����C�bU�brV��]	�L��;��,G@��r���L׾��<��P�=���K,�&jq��Y�{q�5���(�6:��{r���z��#9w,����O#��꿟�%��P�*� ����T��B�iR�_����u�@+."�:I [�C��.]
��N���������"�J�G�4:��s����͋������|���25k��7���J�F�kr�K�AQ�f<p�Qi~.��ƻ����@���i.A �f^�͞0���&�MY.( �n��F���AO8�/8�=|�e����#��q����B3�Ǻۍ�f�q�<�8��0�y9-�}�b�˒����b2w��o�`~��~j�I�s�d���n�U'�ԓ�*�������ZF4��L+K���i�L߭{{�_ p^��ʯ���8���k�[�>~)ܮ���'�Ɋn� T�����	_|����&W����4�#�w����:�ʯ� ��Y/�h�c��K���V�3*�f}-L�_k<+��:h`>�b�*gRu���o��Y�����df~�?�#rg?��I���
��IMf�w|��0���r�=_-�fE����ř䗃oG``�Tl�_�*��O���-="ބne�C���j���E�������CbG���>���M��Rb)S�����(z���f%�Q���kaA����u��ߺ8��]�L2�n����̳�L)�-�	�,&qP�a����|�)�;�h�&�*�)ۂ+=����<Q�1�,�?�~�c'q����X^\:�!H���߰�������=���e����o2����a^Y�����/J�O龁�p�cvِ��++h���O^��澥86�{9���u��F:]4��{�� ��?��	+<^����v��͉?v>w!Ю��e�P�qX���K���< DFC�'��!"w}��"k�sV��/���<��f�W���jm�p�Y��8n�Ŋ�	 {vC�o��2l`���m�T��I����%x.&���oۿt�� 	�@!YMKjLM�����zjt�*����9;+��Iz_��@���{>*`I)��lC��wj��B�*W	�Jĸ�6bj&ch0����9� |*w��q�oT^��ٓ����%,�G�����3�3IOJ͘!���͈�z�4�zw*N!����wwsv���o��o�[����f�|�N��Y�1��w
�Z&�[76�����]dy0�X���>ns\��f��2>�Ⱦ��>���n�+� ��(^��#�3 �/:�S$h5	���sjR�x����x(J�by�JT�� G��(�J�����f2|�p�J������+75����HFx�U#ܩ|��_д�����j�D<����K�-�S�aS{jT����r�b��SO�>�{k.u���+��t�j�:|l,T���l�q�K�e�U�M ��F���!�N�=�0p_�Y.i)Ẁ��nэf���*�d�w�U]�Π�2�L��R;�I��8�lJ2�����&��*��dYM��xɯ����y�	�l�7^J�v^��ڽ
�=Wy�i��S����� Yb+m��^��Լ��\|<�S�a�S)��;�Bs�X��lKx<vR�������(�&Lq��Nm�꼔��Qv�Ì���<���"\�#�������۠���X�K6�S8{�o��e�\>��ӌ���}���ȓn1�e8���_��&����x�y촺�?�,B�x��_���1�>#tS'��j���^b8b.���Mr�/�=-q�W~ٿ3�D�m�Ge�t�=j�2�cS|}�C�A��1u�h}#��@��Xf�:��j��\����\Q����m�`��!��ȭsu6#����_�b4�-4<�>[E��I��q�C#����wL)!
{l�+#�Fɲx���@��-86sݟe��=��2;S�7�������4\�EϑCǭ�&���?���4vA�2ª����-�S��2z͎	�q:k ��#���Q$�P��mqR�C~�����>��#8���p��wPL!}E�$�\	J߃�]�ƞ@0��c�����a]�Y4��QD ���4�=����b��'��'�V!�V��{*�?��	x�Sߚ���{D͊, ����+rw0AT��Tr?R;f����j,=.׌��J�UӨ���-�iw��sP�K�.��	e�l����}@h�2g�5dN���9WK����';wE��qG�P���;Οy����p�vk��^C�'�q�hn��Ѧ+$�k�=˖=��-XwZ-���侢��0�9��m�`�`볚`kچ�3%E�[vb<�����`�+nPKn�X̪�F*I+��?�rY!YE�k�b�\h��k��ع*�@�Z��R�Y�x�~���u�n�?fM�b5��v	o�ox{"��/f:�C<�q��ɘ[��7r�A8qD�Ӌ����uP% �	����g,l�t,�K��f��:ޝ������f<�[�e�ͅ^*"J�M육�8b�U	'���+5W!�fQ��^�B;�ؐ`m*ںCT��poPI���s�pOpc]�ʳ�-8R��qҦa�h���6� d��Sح���U���:S��l����_�ҳ%�s�d�������a.�Kƙ_)� c����W�1��Sa�3�p��W�9]�q�dн��H�0�!.[镍�)C�4{8p|C�r@	�Z�/$�:V/����?����+u��Cb�>i��������tω�xhV,����8������|��� Q:�8��9h���Y�n_'�R�BǓ�.()�a(��oTo+�u���C'���iHe��^��R`���>+լ���)�f�Ұ��\3	��v���N͊��OD7����������p '�j%4�(h��gt�@{������#J��D�>c��r$ⱔ4�G�2�y�M�R�[�=I;G�C���}ۮR|�����tX侬�g�Ϛ��3���Ono�S�/$�}r����Lk㦚�W��ϙ,��^.�'�Q�#��)KW$��,��1�����d0�٨��}"��H,3�J��,�k]� Z�%�l&���T\�}#D�S�6D��	MZ�Kr��1�rA| o���2�@3hXT�o����z����a-��>�$_�`M�?��W��F��]��D��A!�9��L�!EN�z��3��b �dv�6}�_:w�D��������{2�G���z�.�`���Ь���v"��G2�ejHT=��4���n<PH����빝�S���0�?��y�E:?��	P�r�;��3�@v4H��X�s����F`�X{/"{3r����]�D5�P�s���na&ז�9��?*.+�|S/��X�k@D�l�=V~ɡ6��e�M��ɣ��)���t���#CIOU~0G\, ����
���^w��NJEUW���h�)���C�r��ӽ�Q� r"�]���{Eq!�O�D������]�C@���Tq�*�3�V�~C~E��GlʇV�M�bA���t�1Jp���x|���1F�ߍn亯�mA����JN�xh���ۧ.�����܂Yܚ״q�L?$L�g3Y}iU��te@	A;�m�)9���\t��R"�_R��p:F�i�F�EЁ��]l`X�9��u��1�'5j\K6}WwI��9{����@7��t���y�P$�3�?W�)���%��-z5���
�l.<&&��ϳ�H4Vu��<$�f��x�ZW���ZRB�$���p�}!��s����LG�4��W���Ie3�&ԛ��G	ׅ7��x<�|X0�K�C��N���
���4ǖ��u�����I� �`�x�#h��8�j��J��DR���05�b��;�212
������ݓ\#)��p�cT�u(�^��ɷv!5�+'�����c�oP+��W���6�R�F��H1�\�V�V`���>��&�Z��>���M�H$7�'�q�{`A����,�lg�d��+�[�s_�&mn�4䬋���x6��h�Ҟ�>�?����*-����d�ˎ!c|ڢ���w��ca遠��F�D��)߻x�"Ο"����V~������z��w�2�m#�@*:�T�&�����F��������݁��MN�%�d3Ɖ5e̞S�}g��1W�r�Ƕ���z��h�
#�dd�r3�9(����pr^[��x ����Hp�$��3�ݮ��H��t�H>��{�Y7�!;UbL�-�!���RϦ���|d�\�M՘�i��O����"1B�ĲE�g��a��g�����{(]���u6#��,Y��$�������͢��/��]cn���"��;��W�o[��+��(g&[��'exm�-����i�{���� ]�1~Ol��؇=���_c�'CVR|����X���H͐}�����r����VC��T�G��^�-M�kz���ܡ����O.z*th�j�;C��9���_��׶L� �2����S��g	;����B���1�:���?4.�ǖ"�M;|�+D)|��!Dn���ӈ��r�������1�R�a�v'ur�J5s-�`��>N�@su��r��b�z�Fq{�.E��J��A��S�@�G*� �P�F�[���G[�څ�9��Y����T��@��pt�^�)V�S��Jd�.	�#���k��P�Gq�
��u��roUd��v�}��&����'��-7��y\WU4�k�b�o�1*ذ�x_1厌r�w|�B�O)���2�]`��v�u�Tڭ<����#�SI	�s�~=�<2��1��`�^�;��8mO��h5�w'�,K�K���x^�
��O��jPpS���q��EZ��uf�cVv7�H�?��Zc.��sc���̓��'(�t	�f�߮
�`||�､��g���H v�+���U�1Q�볝�u�,v.y���.D��~��t�7�DD��e��a�6 f�^���@�}�RUG��P� �4TmO.15^K�9�Ri48�����5�mu{���m�_�֟�ұH�$���*�xS_���0�A�X�G���<P�.
:��'x%_��%D�X�;��w�n�e��fF�}�Ҕ���k'��*������A�59�Kx!�Zh�9��>&RH�jqy�+�c�	%�$'��s����p����R0��U�����m����r��}`��4Q�#f�] ��U�0X��z�1���ݱ8G�$������V�g��gbs�f����~Z�<���+fa��	UwX᣼]��,��ێ8%���G�qm'�?�h
�C~���+i�9I�����ߡ�}%�����Ʀ}�\�=��_M,(�'G�D9m�⫠�ws\	Q�e���=��w���BH�O;���9n|�r��]Ey����o��#h�27G(�t��7;dkf���ʪ�yT���+0عP;Y����֤!㢀����z�aE��L��_�( ]�^����ˤ�o"큟bE3�{�EY� �=u����w|�Q��W@KF�'��-������I�C�~��#(&�U���7��@�ⴜ�V�C�����;�ڈ�C,gpߝ��?�IN�q�J��-?�u��Ө<B����2c�*�Q�����9�٤�L�Bfq d\��z����W�UF���Q�R��0٬b��6A�����UZ�[�J��S��M�q4����G
���X4�}���E�@%�Q�j@�T��00Q+C������p����������5��2C{�N�Q{D����mfG�I�9��!F-^UZ�j���~e���V�Ԟ�a4^w��.l�)+�#1��*n�C�a�������
�G�;z�w�g�)�0� q&O&X�d����L롿��I��4��Z���nG413/NmT�A� p {��y�i��g8%��;}� �-t�>����|{0��{df�iĳO�.&�+��C,���E��^\��ix !�D�$7W9�]��ڬ��Y'�b;[������Nl�ȫo6���)4<��g3���[��Z�߱mZb��nLu��+Aa�=ơ�\� S�
g�� ��������L�	�{B�����D�*2p��:�T��������C̑�7F�]= �.�v�`�?�v�
�O
z��^t�_iWl��ux�b�'"Қ�'(���4����}"�n�Ly�Z�v����W0DKP��Q9��?y@bV��|rӽ �����b��}�*E�?�U���  R�	����I�r}���PHj�!R� �|1�B�y�(T��ʪ�z�6j�wz�vg2f��#�J��gn�,ϋ�~�ep��Z��ч6���_��[Z�
C�j L���%y�J�l��z~~]��D�M�t�
�U�0L`�s�8[Y5TtHļ��k>���P�x:��鍭��~�;�Y��u7�l�?��l����MZ�`Av*����=��C5,��t�:�TmvA�]I�I�	�]Vav �w|�6�5-�,�$��`�h}��fL�L��#M@�<��V v(0�-m���$K��b~���4�������[��|D�F�wɋJ��Hvأ��-�#�2-��ɗ�7�^.�"��VLO0�\"��k���cz���#D/%JTM����;Q��ڮ�7���_re-���y(�����(�Z�sn��_p�B���D�ңS�/q1Q�4�Ό��i�:p�-ǜ�-[�6�����4R���jLw�_�d�Pj,� t;���A���T@N��߬nZo�HnӮ5k0�Ц7��`��
K7�\���2�1����B4� ��jt8xH�ו�����,�_�&eK���엝gQ�d��k���Ha��h�Ưu�r�gߟ��nͦ�LԌg��7>��'�W�
�*�a�m;���󟐫������~wh���.��k�ז�mL��v?VmQ�>4�������ơj|$.�_Ԛ�'�pL:�r^}~��d!����r��v����mNV\B�Se���3�35E;�Kiɡ�'t��Lj��B,��K��JGҠ�����W�H�_� W�"�.���/��}���&��Q���D�Z
-�2o�+]�ي�tX{��~D�0��q�n�F5":L$�>&W�My��yL�ے���O�ȓ��5��8!�C`���Xsje������8�xp�$�R}9���T^�������˚��EI���\c@Hhr�8�ONB��*'���lb��a���`J�w��%mpf�ӵ�g�J>'�ȕ�4�(W���M�5��i�q����3���6��7d�ri�q/ɑ�6�`��I�,����=ႰG�[$��3,�̾�i���eyy�Q@�����5�S�gï�r�Kr����(,ڌ���O~���bh~�(�CY�ߒ��P$8 �����U*��gQ���o�\����<RH��$��U�S=��Tt�=|b���K3�f0���Vo`*%�qЊ��(BJ��<����~œ4L	��KO�¸,K 	{nȂ�ty>����о0�g�X|�e���dG��[�b����Z��(�2�YY��F
��O^YN����z�
>���Jfg��������U@�a?W��'��i������,��֞�] �Wnb�(�GIY�Z����*G�u�c�>~�9��*g�'F��e��?�E�ꊔ���}s��@�bȖ~�@N��/��n�+����$թ��#�/y����vuU�G�\�D�-+��118�~�0{.[��v/e�~*bΫ�����+�h�ƽ��)�DRBt�2�[��3�^â�w,��%#��#���3))c&b��,zbR-��o� X���X�զ���0t�ˤ��IH�B�#S8�mO��Qv���k���M+f�=����;/����n������P#�(k+>�48k������	U�M��p�]��̽�Y�B��a枰l��_�N�h�_zc�T�{'��p0
�n�8{���._��[�U�'Ǩ���x�����s<vx�����6�	�9�:s% �"���S��\�>�
MHhZ�x�v4�Yij�cgBH{']5H���}��NI��/)ȯ���i�RWE���%.H9�]��
�H�3D$@�wK��D��o'��^��ȸh���0�J�"�]滺)(���Kq5�b�~��K�|	��\ra2�N�`;�?-�WX�0��!����e���9ĝc�B�\*j�E�f�dN�������e�Bޣ��Ӥ�0Kή[v��~�Oz��<��ʥN��¯ \�u��9�u\�M⩷�}�����Nf5|�ȧ. N��C���(����@���V6��\��O���VP�@��bz�m6�M��Du:�`v.��jR��~��>^�X^m?���֕����'��α��� z�:.E�[E�S+<&��wR�Dᦿ�����^�k�~��&@�󷡾Ы�0�g�o	g\m����op��k���(�Ӳ����P���ɂ�im��"���Y��'d'�e�Y�s����v�>@S$���P�[!"��/����s4��  C(E�uK�.{���Z�wh�ت�y�y���K̅(�J��%9�tI���L��˩�EG'L
��ȉUQ ��w7g��[߽�Y��� ɵ�n�ϱ��搰�����XWw+�C�jr���_� Z��o^�z���.�6��oj7��`�p8�� �l�"~��;��I,U�5�l����u�Zg'���e��2g��
�%��Ċ�- �^�֑M�P��5�숗K��NM���et\�3�� �pܦENʏ���jі���-]�	Q?��L�G�1s�(�n���u��2��\57�.�p�M6%C5Ķ&O�
�rSz�$�m���*{�����FW��ej�gx@:���&b��yR��s�㴤޵��n|u���C���v���FK�� ����E�$�+5� ~�Q��p��{1_<�P��V����vw��ɤ��חr�����i���{L^%��{׊/8{rÇ)*���R/�AJQK`k�f�1��5>F��\��[ș���3QT>2�AYE�-�I��30L��??7U��*A^ח�p	S�4#�E~7�Q��P���RX?��i�[!s���Yc��6]�#�W�u i��Ƃb�m/'Y�k�4��[e�5X�X0+��<�F-7Jq���ue�|��,m
@{{���d�L5�J��:��#�y�k~J9��čDx���?缀�sx�<�s�A_��GM$]켍\����V�5�F&/���;���Y �C�x�Yjk���y�\*�L����G;���3���5m�0�R�2��_�Β�{T����>;�~�Z��}�����G�+��j�&C�y՛��I��%��~#���)�)���4ܫ�@۠<x��o��C1`c�D�!��2�*��/9$�~�'r��6�?�ΘsGV8���-������!+�i��̱^[q�m�=�tA�;AI�P7n�І��*��]���q�0f<��?���|s�o��Xӊ�?/q5�/�bW�N��������c�<�? m����@�U��"�#���~o0J+R/�D`ܳ�;ȉ�+9�iRa�6ҶQ�*K2_�6W�8.ѡY7̽٣O*];�R*2��� ��$z]/)BY�t�s_{��Ob�W�{�3�TBٍ�m��:s�$�Єh�D�>RI�6�n��2�<x�H�z�S�C.E��w�����f�^n�g�l�6/�w�<�-���mT�3*��`e9Q�T����N��ө.F&�_���8C�U�� ��^��� yg���8\C)ތ��7�o6�\�/$6K|��j&�^��ًD�OND�$Ө�AO�I��Ȕ51�$YӒ�^�	�>�B�[��t�e���M&�z&��@��zFgW˩=E*��g�L��	�?\A�:q={�CqiI��0!����t�������kQrn@h���%bIܔt�S�nL�k�m\� í���~;~�r0�����}���%��D�ñ�9b�*����:m�X�b�F�΃װ �1S�G6���ά8��:}�Yd��Qu;Wt�6J����bV��|p�׷����
���l������ฆ�g(�̠b?t$՗��0�#W�_2�A��|������of���+ӱ�5Ђz���w!��f/\X�#�1� �Ɂ���|�>VRϚ��o�D �ՁD�W��7��h��u�\�T�/�z��2��<[^u�+I� y=e��yr�F%�Z`��k	mM�bk,�O�Mw�.���߶�-Z�T�\p��8�~�'����ނoF[ܬsy�;�y������Q�F�?�|�"ə)���-���}�f�����>���Ȃ~�755����rm�+��)��3I��r��CYTI'�LV��c�
�܊I���~Ӻ��|˄ʖ "����F��U~�Y,���)�'��_���C:�
|�G��;����{��J�U^�y�6�'�����|�N��!�g@�b���6§��E���D��b)o�����2,�0�,����f�f<U�cxEڮ˜D��/���S�C�V�D�~�?�ɫAB��*�	�hUbK�Bԓ(g�%8 �q	��]���kh�?:�0=�i[L�eqxQ�pwl�{9	�IN���s�ü��hb�W�/斝�	f5͌����0����/y����Ĝ��E�4D8P��v�/Y	e݊�A�M������{S�5J|�'</b����|W�-���Tp:)�����?\�;F��T�%b���$��X��6�+�AS'�d/1�ug8�������?ġj��^��ЕJq��.�K����*�V2�/����ъ�p���X^�cr
����x�����s������6�-�0��Y6�j��O�΂ne^��O�dd$9�8Sd��Q�T����}�Ų�����Q<���'�`��g�bh99��=]H��'Q�+�tgf��`߷��i�v{��3���}^�|a�I�t#4Z�xkV���fj��<�4���e�5�S�y� �����	�|a�S����-ո8��ѫ#[g��������h�L,�c�;Q�#�}4?�U�	�E-�k��鋋��P��p܍�fм�<S�ce��r��J��Ј61/��� �����gО{E�)G�7Cڢ�7���*����pu�C3�Rq|+�X�g��|��q�ztNj!���w�.��v�S��Uj���o�R@'b�@@�!��(�?�ݦln|A�)ϝ�=���ޝ�V��2�����F <:Cq��:tU&\&�(�)d�!Y�� �~��=x�ҕ���<�!'���}@j�@��AA,�d)H��ڹ�D<��Y��d��P�a�e����U)pK$h1k�b0��.��[-*+�z���@(ݽ�$S�uІ�{�f��{�"(7��TM��M��xJ�C��VZ<-�'���Ǵ�b��O�����ķ��� �bvMr�	;n�|��4@˸x�8�,Rir��L�S�:���,���J��@�e��`_ﴁ��G\Y>�(�d��f����'��
�hc~�i��8U������S��7<�p_�$�¾�G7���V����2htx�n-p�m�jqW�3��h>�-!'y�q<e ƴ�p�e���P�U��IV����Bb^2�4
����m-�Eq��k/SA�.3��g1�z1 0{L
�3�b|�)f����&�M7?�m�7Z'#��
��T͵�f+T�^a��.Ci��A��!'�O�K�}~ ��uZ*l���QV2�)�`F(]�մ���`�I��{���3���9YAb���1?�+�F
���t�K�Lڛؿ���ޘ�8�?��
[C��c!Ӽ
x.���e����B�)��"�R�����18@Cn�DGXt�:�Y�OJ���?4�"���fPba'�������� ��}^���?5>ذ�`���{����3����{m"�����ϻ����9S��,���'�X �d��3�h�o<T
�E��XP����)�F�D%�SϰX����_����ع�@�#��M�?6��p��V��xu�-#�qu�}���ڏ�^/�w
Y�r���L��I)���q�v���g4I�=S8B�&�8�JZ��kHŦ��y�E�2Ip�ܮv����#Z��틃�=G�Y���DU�T����T�ɖ^�a��G�1T���#j�Lܲ��R뾎���"��Mخ3������k @j|���-��{�߾l.Д��5߿���>�Lq���E6��J�ȿC
-u-�\g��>L19^�c�y�ŢLC�1�2e����MOk�On	I�"`���X��RBja�so�4nҕ>Ͱ�h7�w�
�(�ؿ��S|a�� h��
�o��F� hG\�CC��u8ݾCcJ��Q��j	gd�9�� d{�y�w17�j�V�o��7��)�~�X�g�ƫ~#M^��,�����q0��-q&�}ZL�dBc\�I㾯�\��:yS}�=�a3p��܉P,^��S���9�4ɖ��tcH�c9����E�c?� {i�b^����'u����D!�y����r�X���WZ�������$,�� G���c�l�)��lu2k�c�txYH$�����ʮ�܇s�ނ�T���c*|7}]bBп�����-ܯ�E�H����Q/>�m��*f�pw��R¬���`�}��Fi�D�#�����'�%�7x�eER��N6ъ�O��۔m�<�ƛ���(��n��0���;SUm�8'�+���k;��_E�HdZ���Y���B%61�+Y�|�4�ż�"ҵz$-]@cO��:V�s��]�uD�!e�I���#D����pV_�*'?1��	�b�nMoЦ�̷�;,���\�);F�1��[1��������Z`f��^�ۺ��G�#�!�e'4�s���,ꜚ��d������I~Y�	�z�Eb<՘�ZE�T(V�Bb��;��!T�P{����Q��%��%Q��)W�1��i�����@S�D�����(���I�B'!q&(E�'��{��dف�|�Q�x�!�*����\��1����m�z�]݌٨l��Ϸ"��+���3��\�&�gNg��n���\�D�q>Wg���
��
�O�x��Q�=F�K��D缐!��-��K��Yf�%����W0���J���#�q��$��V��"a+vTy���G�4��G96'��Vǋ`�v��CA��-�6�=�&!���D7h�_�-����i�<N�t�T
7��*r�S�G��P|k)����qa\.����~.�r�I�P�3��}^�_R &lr� �H~
����n1���SRg_PG�,<T �X&�'� ڼc.I"����X/�԰��]ɀfjz+՘�hw݁�0cp?QƢ�j=�=�g,cE�C$���}/��g�GL�Wx��;&=�ޏ$��[��i���f�q��J�D���o���'�.�g �1[��"���Sk�g�'��,��V��Xd��k��^ n.�ح����V߷�7��Q��Sj6�}G�BR^�/|�T���e
6RI����l��������$=�R���RCי	5�xŦ!���v����i�V4��'7A��Gژ���� �//"��{M�v�J�J�g�η}ďb<����B�րP�s*�Ԅ������ns�P�:��\�w�3J���/���&��'W�k=������6q��J��ۇ�-ű��^Z��%�9/s� �bU�-w�.�g��:^�Q�_�;��ƼU.���GeH�E�UJ"ԩa�%l�r���e���3_�#3e����Ӆ�މ��W��b���t�X�6_C_��A
��QƋ��$�f�])��U��*m��ق����c�<����=�5ڢ�hH_��8P�*FG&����@-��V��W)��7B���3�#?����	0Gl�S9yI#�U�?����[tӧ��r1R�,B�A�Q���41�r�a�7�lη�^��:�.�4��?l-�r��A�8�[�����^Y�ۈ����݇��
�jI�S��P�$��q�O/#��d�6oM���k�I���&K]v�]��ǂ�B0����/!U+�[��E�E+3���Ivi%ӔQ��rd�~�~�Zɜ�D�D�S#��y�������r8�K�p2�ْ#���l�4���
��={� O�Jz�ZGB���z���ܹ'NWC�=!��ӎ�]j��mJzDgo�� pZ��@i��@���e�^`c2�*B4
R�g��}�*m�Q�\J�)�ST�ba��?Aj]���_/+�o�6:�2��?f�6��T�A;��37(���rt&�����j<�t���Rۘ��g8��J�$�'�0�:؋g���se`�O���eT]�R@^�6H(�2����M���j�9 ��頫||�Y�"�3�v+@Z��'�&J�j�'�� �����/f(�$o�^�픬9I 1��F���/C�+h O�� ����Ez�T�]aY3͑�Ax���g���(HRO��;����E99-��%�Qq
?�Vf��)��-{�,,I�e?6��_*�|DKpo#Ĝ��|bGP%�(��qaŢ9��n(�84��>o���Ȉ�p���.C-2Mә��V��3��*����W%�ǝ���إ:e�!�M�%���ܻo�W]������[��掊�B������v��e�#�K:+����C wm��1.��m�h��8���!In�$�~Z�c�8
�?�,��!���k�!��n|�׫IO���	��u�rQ���dtv3���B8�>t䴮K�U�ސ�F�@E�T�}�-n9o��>[�"���J�g0����=7B}NUV�pኤ����o���ύ`Ǿ7u�*�Ռ�$�m%:vp�}�0Y�l7���� 11<�AHU��is.�.�fu�4�ug$jB�ڴmJ<Dj\�W7YE>�EtU���cߑD�ĥ�cE��B�pa媭�4��7�"�	��G S+5	�]z>M75/P���zZk�e#���YS�D�B����4���"�C��Pa{���](B5(���}���=PPH�vZ��C;jsp>��V4K�W�#*(v-@������QD�͐Q�mZ�m�Ix�[z�?�����C���_�^̣-�n�tY��p� tJ�֩�@��TF���@4��U,���-�sEXP�g�*�B��$'�2�����#D<��*t��ע���G�` ?�jAq��sPwX]bE��V!�/� q�S���s#���f�S�V�����Ɯ]
͖�`�| N����r0�K�	�.?����p�e{� ֳ~$�`%t��֚]��:]M�P����bh��.�(��!^d,OoC�/<����)�jkU��aeD�]եed���0�!��.��UR�h`b�$;��E��ʍh
Pn���x�)4]|�,�cX��R`A��w�D1=<��I�6�SX`}��u�KuT�ę^�qթ���)���E2	�Y�G��f�5}Q��x(���8����l �~G}����H�?�����k�x�<q���c��L����h2#�!�U�*�_	�|�������ڤL4��^WA���`łV�&M�9
�l�yoC��}�pR����${��d����RcO/�`p���#����� ��S�B�����Q�c�$��nͯi1�єI?7s�ɩ�VD���&9S-�j�4����"�'~'��׭w�X��jӴ�}�%;�HC�M�H��	��W��0�o��j�T�| w[���M�&���/]b�����0T���#/�[�,+����>֜9ҏuY
���أmY|s��ֿ�WI+��pU�2
!cg��݇;�&�q�Ie�w�I��P�^�Q������Ӵ��MHYw���^6{�a9���*J�1���T���ТS*nc���(���`�����g�RtF��2b+���UP�&��Y�W�R}ėN��C���#:�0�o����k}���I�D�=��T���[�e˹��+�������=��gm��]��(}-,JzB�`�䰂�H�u��F2��j;eX64T(KI��hSx�Qע9��#��k�{���)�}�
�,�M���~�]-��E����E�����n$�7��k/Y+*����=õ1�B�Rϑ�M�t��
����~�H�ڑ�K��h�!�4�h; I�t��M#��Ϫ ��l� ��*�a��ܽAz?~�y��m��w/���\�/����g@���a�����*$���2�.��B�M�ɧ�A��ࡒ���
�^���>;G���>D��*�7�~0?�&U��-*�C���QBGe(���<�..�'>��a�k�Y�-&�و�Ά��D�_u�y0 u�v(� �jv4����3E.E̮@��˵]�A��aAc�1	��D��ܻ2�&��$h�ܡDd����2�D\���C�y�����	o�Ǹ�I��̔��cr
T �k�y�p��D���M5�?
�*a�8lEm����_��ܱ� ?�/ώ��?|�,\:Wq'1�9�_�ɍm	_.�>g�?���\P�{���ɣ����ۇHGA4�x��',O�:�//��a�P� ��ȅ�+`�,x�L�,-O�#rB�.��Ƈ�g���;?�o�K��B	(��|b�)Z���=�`6c��ޔK?��5_�u���˒F5moS1��M�ʾX$HD�dP�81��/N��e��k7CY�QUǐO._�����������wA�v�ܵnu��� e��PIP,:���r2�)�X�$F,V��Zt�n�u"�����v?v EQ��W����M�?����i8L��	]5��4���3��	Uп��0�z8@ᔊ��q�{#���ƚp�� �bAi�pgq�-��N=�nG�c�����9`� s쌒~t�RWL�m�EU�JY0v��Ѐ�|T��+`A˄�LH�"���c<��6Ow{��Ai;5�]�ƪ�C�k�(г��b��)wbӻ�ګ+d�i�\l���	)�A�ݩh y��Y���=H��k*,�$E���x3�`F���#�X�]��暍�����H˵'�qA;5yhA�A�r󋀝�a�C�6��C�+k�[@Sf�2��j��g%(���޳�ꉄ�@jl�:�K����YV3~�԰Tԭ�D����es����q�S0�Ju�����w�YP_�x.zHم9��8���6X7_Q��\˪�1yk��]��DV�v�GdR��91������v�/��δ|�I�C�F>�|�Z���&u��s�a/��`��~���R�7�@'}Q�P©���p*��.ͳ2=�u<hѯXA�-j��c�\8;=ٓ��	��J��)�Xz� Y���H��=F���%��lř��pa���%]2����m��ּ�͙���B�Li8�zx��U�p]�@���Ͼ۹1.��*1��@���:%�¬���d��ogy)L�3$+����D���tt����bYq5+�����d׺Adw}�Rg�'�Tkw[!c'-Y��r/r=�E�'C!7SoLy��D�xϋBͽ�yh�|�SY��@ԅMVz[i왲f(�y>�r�J�ߤgz���4k�z�����K@�$�������E���s}�"����U���jG�>�6 �)�s��_�%>;V�X|�����f�|�����mpgo8 ����nRЛ�	�̕�o2�^ �x���?�L\F��|
�I-�d�"b]M !4��h�ר�*�>�%NB��y�����D�������0�%���M�zF�#M �V�"$���զ-�q�N�C��'��[��c�$��*�0�R��5�-�ݔzȰ��@���/!��LsB?K��v��Ȏؼ)�3��v@��ٽ0���r|B;d{�隚���L��w{)�KN���n�\>�k�k�_A��T�2����h�[-؂��0��G11�t�������
����k����/��1��(�J��+�,��_�d	i�x�AU�1�p�B��@�O���~
~�b�x��R��ܼ�ɾE�4����N���FO�>G��0sO��f����i�
42;hx��N�����}�0�	Дǀ�F����}B��p�t��Koʨj���aoj��XI	l��r�'�樣r�d$Ïj���ف�Q�wX��B��6���7P��4�v�m,աμ��f�y����M���k���m�%��n�]��Qh�ZY�/�)��f�S.�*G���~Z	Z{��$Y����ℎ=�c���b%7s�;�L�����b�����r��+�^��uI��B{91R&OZiV�z!���kM�W
x(��	�I�5*��y��+e�%�LI2�W�Tk{\y�gi��V +�μ���%�ɚi�"y7���ñmm���-CI������դ"�2*$g��yz�^�;xV�������G"v�}' b�G~A�^_NUt(�
��s�d��t@��Bm�DQj?���^.�<�U�}�"����o��+7Ǖ�p��&�#�u���!̞�Q�ͰO �OegvF�iEz�����D��a�[{���I�tz웇Ӡ��L�8M��i��݌/*��
m|��J�<#t����Z8	~�̢��T����������&M=׈��C�㠬�Q('�C~n��(�3��0��uI*���dQ�Ӏ*�-�V�#

�=�e��Z��[�AG ?�3w��n'����yq��B���0o�->�7���x3��qk0V�4��2"����ɊG% ��P�is��r{~5r����C�Ӷ�P;�L�u�E�a�^�\/U��!Knػ������h� Ƃmo��D�c����e�/]�h�v|���f-{�U���|�m�)�Զ��Wﴄ�+�NX�������A ��u4�^Cdi%sy���6jGq�>xٖ�>��[ج;�7<nܝHPf4�o��*�L���S<A:�2�P�]aQ:C��j�<���W�~_i+�#�/�kf�K�<�Z���D�{�m�4�^rc6?#MG�a'y�n��?�,��n�88U����gX6)w��,�+-'��1���+�C��Ec�l����?�F��$;�ĲZ}[XŬ�k32Dfgʕ^\�^�*�0�Ⱥj�
a�H���Ag����n�sB���e#S>��?�k$���$�&�5��P�M����#������&JGTo��X\�t����p8l�5�ߴ�4{!Xǌn���|��
�! ���j��
Z~5^�J_+��N6 ���P
0�>�4ev�����ȑ�ƨ�@)�e*��$������Cᓱ�Hx�.�$X�d}��\�h�ln�P�5����}+i��1(�)d�dP��cb��ƯjO�{���;�/�&�n�6�a�e�!���_�h �5�󰲒۱�0����7AɗЇ˯S�o�����`����'Z�>7�5��ߗ�n���C�z�KGs���)ʐTl2����(0�����5ؘ�/?E�=m���}�Ξ�b+���b��*K0�g��A$b6Y���M��R"��F���7�kkj���$�I/�d�X(�_L$'�g$U��2�*Yo :� _�lX˞�&�H�+�N[{�h���4�I��	�$��>[C7TǨ� �K��!��*̆0�E>��Ǖ ��r�Ќr+�RFΆ�(��w���x�*�!S�j2��!��dk�]˅�[�������Ψ������B�L�K��l��ܭu�_�4Lq���_+ĥȚK]�5s#D_g���g��;T[3�u��z�]���F.��S!|�>��11:M�����$Sףc瀗D$6��TcM1)��5�g퓃<악!�}�+�y��b������ĄZW�&�T����������4�֝]$�)Ujb��qѳ$�)�ڭ����U�?Q!��pWC(D��Fy	�co�zOr"=��	5X�ƭ�l���R���I�1A��u��|¾L�?���y@'�!�Y�����E��ɠ�~H��U&U8�8o���a�5�l�#�!�֭�}ߊ�fZ�DPr'� ���=������$������ĸ�ʂ��$I�Q>T2�5��Ƨ��r��M�,鬒��P�v��U���m��ݜKt�*�!P�}�Q�\��ks�̹tZ�f����:�6w�tM�SB\���j��b����@9�߅Uh�)%_U�mމ�r^L�7���]ޱ�Mx����s���J:��.���?�?o=����gc��	���ݫ�Ay��y���j�_Ü�cA���Ch֌!�"^�W��E׼m���q���St(��6��SX��t�9�L]`�N�-"���ct�����p���|8	����E�閬fV��2c�f�;�j��mހ<е��$S�킡z=dkn���靱�q�]�	�����7ܨ��{������6,5;��DT�P �YNa���7��f�*�շk����f�+���4	�����R;ZB�GC��z���1RB�"4m�"q��m� �9t��r���J�N��W����,���}�ӣ�j��5�y��~I+��9�r��T0��h������E�����́kn��<ȣ�T��NW���퀥��&f�ܔ��b�ұ�ꋭ�{��Q6f3��G�ivfM�i	�y��Wҥ�ܐx/54'r��#G]�]�ys1�X:�'Q��jfBX��ZpѬ[�k�8@/wih޸&��u�4� �D孃�l'!NZ&4�Rެjdt*qz~�;y�]U��V�6>������H��'��~�
F��疽���@�T��p��?��@|��5�#���؎KW��%\��*Jҁ	!�S��A���𭱩��,~ͤ�b���G�4>��|���|����(ǋuƹ׀J-�`�g�Ԯ\oXG�Pe�cm@��<� �gK�3��m"3<���Y�&�Jk��vl�[6bX�jY���j�bz���`�*^�0F�ള2K�ԁ�H�h��j@h"�_��sk�7��&:�� ��;&q?Ѥ���a�h���R5�6_o7��������6�i��L�}�,,�r�n��������e���~�������8Sgf�b�Ce�0�n�S"_�A�)����UQ��ճ5r�z�x�5T�ar�ߞ��%����"J$��-����Tu�	���K�Vq�BWa2�ߪ�.+mҘbk��.�,%� ��}*���niD�_-mipݖ��#O�U���>ے;��Y!m�~E^�OI�T��Iu�B�*%����ċ��f��B���_L�*��a��ڱ[G���4�:��_�P����	_Hhn�R����f����.ܦ]"����[s�$�um�\ş��Ŭ�Te��@�����J�3� wؑy-0g!G�S@C��EӢj���V:�RU�����>�O�3#�����[�!��&�/b����Yۣ�J8\�۫wf� �01���6,b��7ح�. /d�0w<��G��z�'���f4/��q��"�uC1�~��!P�=&�6*Z�k'P9Tz6������c �6�K�����Vjs���qk܂�;�M��P�c[�r}�"����]GYx��3��g�s"m�4�l<@���|���������u5�1 
T�a���z�Y�X���t��ݠ|�pVd��d�~��*ŕ-���?M	�K�Z@Y�o�&�����8�D���7,��%�th	��$n���?7}�d|k}�a`��_,G�T��k����B�5��˾�qna|e�Qi�@h����Œ��p���hT��/Ҁ�˜���C$@M��y��f&;���-a����;��?<V �1��	�N��z:Zs��'C�Jd���}�KVH�q�FHX�-������v8�����!]�
�Q��k� 
vG����8H�Pey;�+�R9T)�i�&j�����80H�D��
@qM_Xa#N[��fK����I�Q��g�{����v���+i�1�(���-�+����T�ѽ���"E���VN+6T0Q""�̤޵2!�$y��Y�.t����1Œʆ�^U,��=(���sk�I�phI����sb{��S4��8����}�����j���	�Z[ae ^e���t��K	kx�I�bPF����KM�:A��<�������dP�as�(�.�[�'J�vO�Z��d��,�lsXʞ��1֎�ky��C����x�S�\�������&WӮ�4��ۙ�/A�Z"��{��T�Uz���mpy��s1�y#��Ԇ�������cqZ\�%J@�_,%�:_;���[�*���a�Ê<V10C�����P`P�N-��������ﺃ�F�s26\���^ ����-}&s�b	�^e��컧�H JC�P���	�UL`uM���I�O�\���:j�Li'd*�t�+N��6챥�8�Հ���3����u��V�\?+�.����8:���_��3�T�/�y��FؠD�N��O=�e�8�C�������b�Hj�{��y�����fz��O�_�?<��ו�f���NXZ注zZ��[���v֬� Lر���6yj	D���d9��N�D�,V[�+.�q]Wm8�_����P|D�.F�hQڛ!�`��|T� 鈬P�@������O5A�����1bf+U��8JZ�֘��8��j���c�u,2	���|�&�π�}�9e����^2�q������*�?O�/"Z�l�_�����/X< ��٥b��&�-�ɗ<6;��z������9?|M��mñw����/�[xU�0hwF�z]������禍C��E=�O��k�6\��{�>Srs�Z�<j��mm�[I���t���wM�U����8�a@b��h0�u���P�m�Q?��<)���[�,n��0d'
��	��2��@��i�� �R^��O�]��[��U*�U�5k�Q�h�1���H����>P6����kE-�x#'_��+����P}
� T����D3eO���i��f��H�S�=1�Vc��P�i�I�/u-V�(w��7τ�������9Q�?R�[U~/�Y*���m�m��� 	�#�j~����)�_�0-#}$���~���5&쎲�0?��;sof�ķ���+�����v^�{YJ��a��norL` {�Z�����K��"
�ъmܔ��P�~�͗In�&���l[�FcT�j\�e���&�'SɆ�ƌ�&�6����X�YN{쾕!�/7U�l&�>���t3�ꈊ>��h�-�7���c�Z|=���m�(��{x�( �K[V����������.yxS$H�up~�k�H�i@�R��8PZ@�\�4�:J��<��o�x,����J�@��������>�� #�I	<?@[T�	;���Э���g4�4���G0 QkfG$��Zے�%A�91_3�r�� ;�������ޜ`<�>t���9?'�r���ד)�o�Kxd���=�Ie=L�x�R�Zb�ϯ��%v�\E�Z����/�׸êF�9t�|c�
�k��#{Y�!�������#!!ح��Қ��D���a@*�B���g?��H�q(����O��3_�	�k��(Wx'��=�o.�&�R� �ձ ?ބ����\DF�%RS�~�0�-���9
pj��Ψ��?��%i9m��V��DZu!@V�n���r9�3m�߀ꦖ�;���W�&�^ tc�c&� 1!N�5����r8r�G��g�V/��<����]vw�#��6�L�yȒ�fJ�?�Vt�ώ<�����!�H�������u�C,�`g���*�+���^ٜNmp��p�k[�x��p�x�'ͺc��}NY�� �Qދr��m�b/��AjD~Q���'9�MZ������7;�0) l�Fx��%)�����/o��
�c����<���%�����t��h�'b4��%%^�3�X��5�J�A����ꙮI���С���u@�cުK@j�&�õQ��PZb�"(\�o�͠Î]��"^�;�Xa!�>��ؗ�1@��{:�{�����H:Q���ilv�U��ߵ�����|i�u2m�[@J�'R�؀�җC�9�5�2�9]Mqm�OA�N�Eg��>/�궧 �!ěr�F5n��k[�dˆ���,@`l�W���&��C��=K&PhQ���m }DPu��ؒ�mݚ��JF�7!w����n��#6#�l}?��� ��m`R1��$6)%�"���"��ǰW��z>��K�R��2�W���F����k�=���<,8Ab�I��LG��W0�ȶ����������CHf�=`(gM�g�̚E�Hz^gO�$y�|�PV�_��7vzs��5ԅk������'�_��ll+)�tM
-��\�iKVepJٻ���j-v�s��~>gn�qU̕}�'��$��+�z4���W��\P��#�$�(�*<�Iژ�׮��8��yu����M�]W��z�].◔��8��X�z��M�@���
uk�~B�y2j [*L�p����8:�<o�E�
~�B��ɋ��3�tK`N��8�a�m�*ǴLĽ��v�-�5Z%�軀��C4�-��:�q[d�p�2,�t~I�I��� ՜��J�-�Ym�8O	ۃ��0 <(,(]i�&N��qpc\�V�R��k�<�)����U�K�R�] ��X�r��~� �3�q�B$�8��'K��F}�6�O����V	}��"�w��Ei��\�e�] �ÿ��v`��U�" �~*���� Н�F�p�Ũ��}�/S�M�hL{V���v�a�ԟ��?�\ a�`�x��yo8P(\�nњ�M8��H8B��B�~V:M��¢����an�h+����hM��+Zdf�Йo��]�|����h� 4�����}c A�e���f�x�����[�>J: ����罽7�Y��x�16t�ɴK�o�Y��M�$�f����w���V}B���P���!$��PSc��Y�F�d�=��Hutt�p�p
�.o�����S,����Լs�8�gЫ�� ~�mfK�B4PBÂ��1�o�DAo&��̮�㢺Y[6uDZ��E,�Ĝ�lLiD_��a��L>��9<�ܔ'��: *ڥ{��)H̖��l���:��Q������V:��4�F�{�D�sY'��v�ײ���n�ޚ{���3b/�!a�Ȅ���j]^J�C�g̯t�sZ�%c�V�9�p�?�ُP)1��&�뢆�qHm��4�:pV�����e�;=��4�z��������Е滔ɠ�p�*G����I'N�Cv�Xd��v�9k�Bo�,��\�2�Nz�����D�f&o�Y�#�I��#x�1�k��4�ٻ0�?�E�v�k�W�l��X��^Kn1 ����ic�	�T� T0)���,�Y�s���46y[>��5���c=7%�sfkp���S*�24�_4����k���T��҆��&?AZ� ��]���KZ��#{*�vl)@�**�L&{�Ǖ�R?i(�f+�v,vz���\wi��{���-�Y3�J����m=�
�E%���>�� r�7��Gj���O���<�M�t���3��`ض���i�����g�?4�����nu��1Ѩ��.�z��\�J���|ǉl����GqWb���@OpX�ջ�rӦ#�:�:)�SB��� �둉!�y�,oҾ�7�����k��I�[�����s�oYD�
�ݔk��*Y���D���%l�piy��$�������d�)�5��X���F���V\';v��aԌ��J7[�w����+�`j1�9�J��r�ñWo������[�49�-��q�~kWw\ч7v@<ЕH�Y�h*��^��=�L�� ��{�ą��� Ng!_�}�V�+=.#�W=���7I�KC:[�!%���?{l@t+kq��wC?�D��
��3��H,c����4��&}��:J�f*w����$>c�x�{\�Ir�.Ӻ ������	��I�Q�T���tN��F��Rd���rI����=�I��a��Œ3i�~�
�'�ߍ�j�vAF;ĸ0�=e�ɑ��h��{�x]��j�3%6���>I��4̱�I ���nPa�6n
���`;�	H����J�--�>2���K�3ZO�t����OF`�]R����(_(1��j�5+Aߋu��*cVMM�a׎k+"]+ۈu1-7�!,��]�*眅�{TE��^4A�~��^bb�Y<t�����NJ��Nڇ�� 9J"��Dd�����Ü&�@���e1蝨��ał�!���$CsH�r�$�e�j�NB���\�w1�]�܂���xW�zc{��m~Nk^���F.��Ù�+���Q��{aG�젫'k����]J��:ԫ�!e1j@	h�[�v_u$�u_lȃ�+�s'�n4ƞ&���Mj�ן���V�FR�����mA߅����F5����7U�Wp6�1�G4���0 ؈P$@�@���'�E,�>Fa�(���<d�v��t%�0��?�g��4�����T^����Rba��t�Kl����\�}�����?��+�|�S�\~F`����'_:O;����䦬mm�aj֠���u�'���]-?}�"jЌb��lm+���������m!G]���g����Df�ek�H�Tk�������`���C�2�B��=���8��pR=���g����f\2"G�z��v�P��%*e7	�\"���ٗ~iG�D����܍�^����9:�������� ��f�
�SU�N��d��`��'"�L����%F�4p�K����_`�y�+͙P]��^��ϭ��'���~p�fRn���۽�~�G�		��j�_%�R�x�P6�L�Y�H��٠zzz�e8l]��n�k8g��E��>�r���Y��r���9���7�ɛ$1�LW�8���_�� G����=ܷ���Co6��ȧ�?�����t|�/fB�Y�$��y��pjϦ�&5����h{Q�u�49��zr�٧��/r��:�/�v�I�i�A|���٘��v�.	���JZ�h��i<�c��-�MM�ߏ�ڴ��jc������Vl�^Y�|�z�_�R}ݏ�S�(��1� �e�B�� *o����'�d-�ƃ31�+��~�%�҅D�����Lx#�a`�t
�0u۬������>����r� �:0�d��?6Hy��a�l�C��MR
j1�1�^���~/���W��"w�5P�b}�#�T4h�+��ƽ��FP�PX剂f�b��dʼ[��N��9�Q�'��Gč�)Z\p{c�ڑ{яՒE�������ݍ�. S_Y	�R��;�%4�������n�A�'�����4O[HCۭ��!䙬��(=jwpk�%�\�`��}��Mb۔hUA�W�u��U���x)|rw�41�X�V��3D9��h
�7m:����]_�.�΃f���~�(XZ�j�&YA���w�!�+Y���4��.�4-�ϻ\�M| �P;�Y�*�l<�&��S�����"+rNK��/��jZ�1jj8%��xy�	7�q3�D��u[�{�V���q�����f:g����8�2���Pe��D�T�0�|���G�di0%�n�k�lʣ:��x�"�$'u�
�+�qm���<# ��	�:�=neld���\EA�Ľ�+�u,&PJ�7^����.��� �K���!?eGR}a�G3X�#�T��z��2�m�t8�K�\�'ޣr�UWT���'�6Y%?M�!�z^%**� ��s����p5*���
����2��I<�./�E��#L�W��������Hz����)�a�fX3�mȰ�1{�xz�'�jь�xH���B�7����=�\���\)'_Kr9H�CP�� ��cv�j֍N)��:��XN��j���i�kr�ZaK`$>��ѧ?���X������~S�nO�Z�ũ�)H��a��7��C.����ʭ��	����z�_���$uθ~OQ�ҋ���`F�5C��o܉��!ww�*4�B[-���)�_^'%q���Ʀ��/�՗���A�22���a#�W���$p�}�+ f��N�#���6�<`%���Jz�������]G�a��A(�)�����˸�1I��Ԉz[G������P�����,	��c	/����g���Z}-�]����1cP��n$V�r�>�]�ia���B��^��n�s��!q"��{7尾��I��i�;N�G����񊂸������Qu{��')�����%�\�5���".�]F�3$|�ES��a-&�"q���V�5U�6ae�hIX"
���ǫLw|q��#K>�����CZ�@EAI�:��;>Z�±H���W8����C���*$�%����E��
�#��4�l˞���T���h߁���^��>܆}wf�%�W���\�C���;�]+xtZ��(�U�Ia�A���[���=�{�`+��R���.ʷ:k��6z�6�c�G�D�6�'���~N��(za��b]՟p��ŵ=T,-U�L��`��8�l���!����o�^t�v�S�Ba*���aBH�I�
&+�-DԾո ��i�Q��cja=�{��eP�_܉F��{�Q�����c'3rpJ��ru��)��!���Ri#/�w���S?2�s��5ZN	�!qi���j0�r'[�[.!�'LՅ̝3���8r���n��Kg��C�c6(t��o_D�bP����o�u�_����	O�*i�i����TU�-5�p���v������ֱ��.*�hh�-!�`�%-��ݷU��Cv���������N5c�G�6?~ŻJ�*xY�c��mV�M(eHKK���>l�c��� ﲩ�����Ɠ�Ņ_�=ʤ25l�U{��'��)-���?Z��� M���IQ$��謉�$�'�1� 6��_rm=�	�F���<�4؄
f5ܥ�,��\��p����b��͛P�{LT��Q*�sҨ&�F*%궁�W/
֔����N���G�"=�W��!*֌��c�j�ό�^�Z���x�l�R6`-�gT֢�Bo�iv ������il��n�ȃ-ܡ��`��ʀa:�;�%�\��lF��V���`_��gt_��W��J��gG�/�h�����XH�3�]'��|�l�/y���Sc�'�Zip�5=�i8�U?c�ߞ�p��e;�1�C����\�l�?��/������Wj��d ���?���f�*,�����#��aS�νc���G����.O����r5 X�mV��ϒ��R��8���klF6.n�w��c��;~Kv�ܝ��V�,��y�",�U�,}'>�N����W&�5��v��nD��������O�,�;�E%� ܻ5��j_�4B�d��لm>RC 
�!��[��|����j�?�v��`�8[X��q��3�$kZK9
>Woh{r�1&�xryvԈ���1�$��s�	�?�?��Tt��,+��=���Q�J�&��߉�U ddnطeO磭lVCH���[�\u�e����@*|ؘE�Z+W��:>�B�d?C+�~�3��T �C����xk��BU53YP�Q~"�%��4���U�ޏ�쨐9����T.	���2����7	���wdF�t��n'l�N�꫹	��v�-�.�L��l���B��##��O<�
52��D��b+�p��$!�v���\�a��s��'�vݵ�L�t�x��ȭ�����YQp�I���C�TD� � +]D(��WOQ�ٸ$}Oj
qx�a9s����曤^v@dB@����}��C������"�;�� �~��%ޝwM�<���+��C�+[-��?�!<ɫ0�(s�Ş�Fw���Dg���H�<���ƺFby�6R�e2+{ _���,~bttT���Kmg�á<�Ix�>��t�HBR�(ʹ'�?�6�����Zan<���,�W���XT�(܃=��㲤���������%7 >��$Y	m����.�=�lS�X��j�;Wn��h�꫙�4'%�D��C�f>Y�����	F�){��Zb͕YQ؜2$¨������4�-���N;�3�:��P,���
	�w�jjNˌg&!ZwnF�!�m�y����d���D�#��
$HYvDf�}�y��$A�&^�L=RC�ȁ� u�����ߌ�����SG�)�jT���TY�ID��ۭK7)���A��qE&4Om<� u�Ȥ�k���)�����EZ�b=��l������l�i��;m5����
	_��{����tXd��A/$s{аcA�d�3�^s^7�c��MY�JS*w�C3(���7�*O@�ZP�9	�ł�U1C��]����6����� ��J��e=E9,f*��lȄʵ~bQ�!�%��fq��?W�B���#���������Q��o��&���[�3�����8HU��+{���k|X& j�Y������&ҧJ9X��y��3�|.]
U]/r������o�����A�̣g���D��9/��
�d��]9_��̖�A��=,7qbP�* M��hF�ǘ@g4~��%���j�����|T��OD�|vynIJ`�9������=>0�����u
5�o��\f ��
����d�ܤ��3@��ވ����yN��d���C�:��Z�uB��R8�R2�N��f���3���<tW�I
<��?):�ή�i=�}�eSV���,��~M�#���_���b_J�n��OwM{�S�����6Y�le^@0��&j��㧍�X`�Ħ���]�W�rmO�BX��zZ>m�ARr��0��	�x,��t��%���+H��>��-�g;.�.���4��"0T�S&��L�����n�[4�<g��g$��ls�wQ� �ف^k{�|�9��o���e.?��������R0���!bz.���.��Ÿ�b��ɖqՅ Ms���W`G�?d��������0L3��c��\>[��6q�&RZ�u���	/��t�	�/:�C�tݟ�0ߙ���L׺�ow�+�o�Gz}#}��F�I�#!�u����-�-�a���f��I�Q!�u��(z^T,��������9�C��3�~Y���j���ݳ�͈�:jz@�V��<�K��8'�7n�8��� /ޛ����]p �ZcىG�K�@��w����"����M�J���X���h�so�Z�T_�pՀ�1�A�DMp)9��Fqކ�N�rli<·̩����!r�ϒ�� 
LK�n�ۉ`�,ߡ�/>p��^葃��k,�z3�x�������Y�;�b%�)BS8:yz~��f��&�j�I�J��dd�u��mn��\pLcO�![S�Q\��1-ﺦm�䬧:�?�)=�`����T�>�H�W�	wi,K(
lc
�@#y_�W:�� -�:���AEptϝ@��X���P��2���k�4ȅ)g������
͂q
p�AJ3�.>uв�b���Y�����2�:�k�W��"������9���l�&����X�G���ǻs���kk(� ?�|U��u�U����}����8My��\��`qW���G߼��e�
��g�j�]��nB��O�EZi?����[�� ��,NǬWP����1��2兽Ǔ�m�qӠ��0���VC�5<����s.���3����< ���K�Y�u�4�"a�Be
{�@狄a~�-�截n�f�J�Q a���+�BS�`y��ź��N�w��uY!�R��2l��lDh�K�%��(���A=2��r�T�G�Z���Nf��<!|�n�}*�_(m/���d��k@7X���ቖ$�Yr��=Գjv+���̧��ڹ��6fre_i{?`٢l����jS;9��sZ���r��R��)��m=嚋?�$G!f��I��Ur��֙$knio�$ ���荗!����>�$�4>*G$�F�_��#i�B����۫����Z��N]j:�ۻ��1��������(�RF�2��w�q�d<�f����1��:�:���Z5}�$T$g�}�ܾ7�t�=� u��t���A/��(E@��*K�3�tO<�zf�I���%���2�"a��JJ�k��Pq����".n3*�Ӵ����B�0�����>�^B@Ȣ�'&dχ�U\8�%�21o/jz3��9 ��F
��Q�*e?��j�2~�V����W�z�R��"_Del��#F����f�0L�]�R#}���l����k؜ڛr�VǛ�1�Y]�*���!�3��;Ӑ\�?l`���򢼍Z����i~�(hSoD��3��X[e}�8c�j�Cet���v��Z/ �:�!w�l���KFG�r��AW�һk�˫�SҀ�d|��m����_(0�3�6�v��S墪�>	qt_:�úAW#+�(.ߐM�v���W��<'�&��T=����ÌJ��)f�:I�Ү> �Z��P��p�W��1k엯n ���L�c���qr^�(K.��nK��a��~m��;)u�S�A�Oy���a���M��L(�˚�sH�%�;����ɗr��|J@݆�[�*:S FT��[/r�X�-,W���f�C�.0<Y�x��6@��7�:%^ȹ��j�~m(�'R2��l�vE��G�� ��Z�4ʢ�H�1���=�?��S������z��j�P���ީ���#�3J�O�*��NX�Yѧ���w0D�����=7�|�������𕘦n��V��e��� e˨������92����It~(�3���W,�K����(\�U/E狾�0���i~��s#�+PP�!��Bms�i��1f
�;J���:���M݉@��&�4��"�0�_`4���� G�P�8N��] ��m?�H<cvL��W����ہ��~Y�C�-�m�_-�5�R����d6i���ePa�Jy�_�צޚ���x��+/Hb8J=���
��WP2R�߈'�֡�/���1�h�bj譿mӘ
�@�=e��˾�9�bq��y��;��cF�@��ؚ=9�v�5��/�Ҝî�6W��'x,�N@Cfջ))Z���F�,�Q���oW�J:R(V���<r5*��H!I��'Bh�!DMn|�f��tsi�q=�n:�ԘcE��P_��J�d���}Z^��fnܸ��⭂S�8^�6�c��j:꜕�uy*�ΉO�F3w~�<����_=�u�`kl�x'gn�_]0���Q�& ��zr�q�9S:DG�Np�i�����)p�W�A|�X
����Ķ��q=�sI�,�j�է#�����H.	��Y���/��@�\���6��p�a��
�j���b��7�9,'|����=:L���,cp$�^����na�L%��誅�/�
�C&:�=�G־�Jxf�7�y��V�i�dgA g�޻�SIm�}F�z>&nCa����:�e����ԑl[�b����z��<��!Y!6ߋn;x��9���3�bN�^����t��PM�]��1� rݪ����`N��x �+g1�n�Bc6��~&a�����S9A�.`�������+����H�#���avc�ﾟ7�/�P���F�ϼ�G3��8��y�
nm0n,����`��zci��&b6�)�ҹ��Rj�	xEo�k
���r�R�qۈ���܊��	�F�1,@Z�ƥ5���P����I��n�͋�L	R�spK��ٗ���Z,:�}��5.s2r�`f�����!z~�����HZ��!��n���k��3���m�}�u��	�!���)2q��Ck�|lA/a2�^�K\�H�D9H�8v|�h�Jj����9	|	�J#D� 1��$Z�,� $��9�x�S�rY��;U��4=
V���
��2�zdEΕV�����|�!���1�qbH�%�U���Р��l�{(c!�Y�\庤*b�<�,B�#=]�{@sny3Ʋó�B0HU���.#���Ǧ�f�䯴Tb����zNx�7+�fT{� T���i�&{�s(��XW���ϵ������x(   ���J=HP^��8��ʟ��Xu��4r����<xZ����mO��Rr��;�~�[�Va1�&���=�Wګ���n�7ؿ��04U<�tg���8��&.5L�J#|W�b=]F[udL9:��!:[�rѾZ����A�6���Ǜ��3�$<�&.��b�(�#�8����G}�YOُ�]7w��+7�޺6ϒD0*I(����(jF�:T�)���?=��i�Gg��e���&�7O�0�m�3��8���<�bƮ��q�U��,L�5��뭂��M������#�����z?�6�nu�w�vgZl��ϱ����Q-�,,����<�WMw
�"������ض(�r�>��+���1'SW���H�����s����dhW�;K��/�!��%q���NT<f���4�`i��#5A�zb�&��M��Lx.�����_'�j�����a�������>_����b"�]R�-��=��,gUn$:�dKeR�N��p	�k�i��l�ι�sg�Oҽg�j�]}�9tGNAA�%L hym��+��Ɋ��5j�*���	ʼ��b������u�������E1�efS�����>�Ĝn-L�R�r�O"mK�`�gеf;F�T}�aᄝR�	��`��W����0�2��$+)L��.���$��&���_X�Ӊi���c�i2��ښ0���h�G�{.�h\���D���V�1�GQ=���{SC!�E�<�%`�K(�*���w��_pЃr�2$��(H�u�U=!�s�K�CK7�a8��=t��<����L�;|�]�с�
p��(�җ�:���Kf3���f�o�����Ke�{H۾�a���'��
�b�"%t�3iiusB��`�y"� �OHY�xU���ט�� ��-'�����,qzGfy��.ﭾ�gyp�_"�$������fo�.zP&'Xw`���4��*�3�d0g[2e2;�,u���̇f��#�̢1h��������Ƅ.lN���WȠN������"DuP�_�j�?��7��ͺ}�<MC֯���p6M��p-D���!�Xt0�$��p�ZA�����i�#����C �Xg��rF%ځ�,���{��w�
��=�z_��l�4�Aƨ�W���v�&� �QBnH�[��
�f�+@"M�m EF��*aY�/\�<�6�������CL{w���0w_~��V�b�f�>Վ��y%�<�|�,�_X7!�G��Cz?�����xM;��W�M19r0�y����
�逍�6l$=�'�[�2�k�a�ޝ�y�nڍ�Z�U��Nw��u�e������g��?Сه>�{�z�`�mX�Q[��N��!^�	�2;(��7�>���Q)%&�j�j��Y&����N\N:o����\
�wø�%�Qr�Ó��7�����sУR}31�]hp��o�/5	t�L�<k���b�8ӹ���ƶHOU�	���׊�Lݓ��
]�<|��u2&3��Sm��:B4�{	�qNݵ���α�$��NN}�"쾎�x�(�7J� o�G_��<���cZo�DDƊ �B�=��z����C��p[_]�L�K\�J���>�;"76|��\��	�e��(/��̯����\����I�?���Y�N�ի�F��x8�#��RpcקCu���z��֛c����cv}�x�qv���4�xg���3�8�?�	�"T����4�� 3��p<�;�ݜ�⊐���F�X��W��蓞��x�����X��v�z��K.i��[�ټ��q�O�~\�ރkA���̢����ع:�Hm�T��� v�1��'#Y;;�yP�iPޱ�aW#.8
���/�������L�Y�lM�A9�ۂ������TgQ7��lZ�mω�������Er�x��AM�*�by�zQ1�)����h�F�:������I�U=�!��h�K��U}V6����X�F�F�&&�)�B��&v��<�(�ǐ*L�Q��ᾫ��z���~y��X�/$��i�צ.0����+!��W-���=��j��Y�B�VH�r�wË���$7�>y�rѥ;�f_X�E*��}�[��^���z���Ő(��ȧ0L�h@���]I�l���o��V�BkJ���r�n�";(�abu������a� �]�I�����<�e�6Y����`#��3Lҿl�&8fff��FB�ͮ�{ b��[�>��g?�=C�����w20���b埒3i�:��E�7wb:� �hi�1.��lDs����{������`փ�s��? [���ۡO�Q-dKQ5�12��P�8iY�7�Z$�xo4�����*P�t')*�:���lq-���|��}�g�ϱ�'%��K�O����ȱ�oJp���6}F�b�ä6b�S��}W��Lg�P۷����芽b^����Ź��d��%����s��Gi�����ծ{�k�Y��J��J����3��HN|=cCvW�QΙ/��y8e��%�"$����X��Ǆo[g�<?��!Q��q6�|�F��ă:��K��Ս<H�_���Ɍ��e��pZN���vT�n�nV��`��uF^��W ��������c A�����Lk��ŅF���[�UU3L\@� ���ʤ"��K���F胙c��~r�>�S���3�]��3��k�2Q�۶�����Nh��2l�|.��lT/c��V�-߫d�:���e�� ?�\������]�m�5�Js˰hJ�3���y�����;>�ӈh�����m�vQr�N�N����|5qu2�CN_ЇV��<�_S��?"��5�j�R~<���4�fnt���OVU'�A=>	�,T�a�PX�V�Hnx���~v�� �dv�h8�炉 T̠{n !� �Y�N�V��5��h��_m]e9/G#��>^j=&��v�����p�� ����]qי�Wh��u���ͤ��QԿ]��륀H���Y���hm��v+���J��&-��hf&c���������x�0�ƞ �N�8�>��W��肷ț/�����S/%L�x��
;���pѐ��������k���2\e,d"l�^�z�*9l�0��M��g� i$�k:��K�wq�T<-r:�����M^��z�Y5פn%-�ɣ�w˾-DҺ�W\t�|�j�}p"�[��4�4UЕ�,�{�T�s��L��
ʉ�Xkt�6�����}�G�����KO�'-�"�v� "���0ʑ��V�"��^H���'�>+I���4T�n��zE[�����K��*���m���?�`�k����N����s�)F ����)S=^%ἓ����;�}�ˌ���D�+��	aUL�n~x��nv _m��Q&�o��S���S���Ё����כ,�ng�^��_�9f@� ��["ƿ��~��1���H�E�1��"��;ɢD�%����e�hՒ,��r��i��{_i����G�}��]3f��q#������g�8O����������l�&�l%�����/�4�����x8�Ŭ�Wݲ���5#/M	�h�_�`ן�jW�CFP�i��=��e#@�C��XB���|��=(�7�g�͛�o�p�����j}oVo���|�A��M�N}0@ګo*�R��p�s��v����x����x�n�O�j��08h��m���fwځ-)d�\ʍ:��F�'�kqm�1Y�fR����_S����),V�E��ω-���\ci���6yw�6��T���Y|�w�	{5?�� �����V'�T��F�\����O�av��y�J��KN]E��A�=5K'p�P��rkM73#��ZUyV'>"����[n{@Ѻ���s~"-��h���r�������b��B��J���^�k9}�	�����l$1�@tN�.�u�b�����4�m�� c:������|��3�˳��z��
3�ܠQCE� $ę��p��{[�3�x���7;e8Z�K�A*	������q���3�� a���M���c+�˴i����� ��k,B)�id�3���z��4�r�쮩�� +[~��pP�^�����;k&�԰��
-b��J+���bg�u�oQ��*Xx~����6&Xhő���=u�!��1��	���Z�V��0F�
>���F@���F~,���g�|ǱR�<�R�e���D
D:y�u�<��mT2lIX@P����՜���_A��`V֌� 8}�� 8���'z�*�m�&��;I����ɖ�W߃0�!�:@Y/��K��P����iz�����/޵;�.b�Y)�F.�(8�\�XR�9>�[��Г����?V�J-w�
f�ʾؙoy$��_��W��A�*gj�Ҫ4 ![TP�a/�6"�B�;;�@l��j�zTS/�~�SE�i��	�l
���ж�mn�ȞMHQ���
�sz�x~�����rYN�ğ>�Ŷ��%H�#������t..�z>��ib�v��N`)���"2����?9�G�թ﹃�v�C*�ºn��`ִd��Cz<`�aUv�������(�|��W����_�}�S8NZM:y�s0�P}s��t7`�V�����d����ͦ���零.W���~?��kI8�9�Y�P�����ٸ>?�xx��̌���_�\h��zhX������t�.
D�2@��7[6��Ლ����qh��O�!D�n���"�_�(&�|a[oZ���y��O 픆૭!���fA"-;w��U�λ`����W��g�4�AC�>t�����O�^l]�+���6�������ѸR#�&˺��t �G?�?��>y��u_���"|�2���H���)�xܢ��L)Z$�����嬈�\k�.������#����_"�����ncO���Y	�
��Y�!4��0����k�Q���׊���HV�m�������⩲,|8�f�mem{�o�<-�HT�&G�ra,������ȁ�Q)���r�wq��Z1ǁ^�5�an9㒑�L ���ozD��F�<̾ߗU��q�N��L��O{���b�1�k���ݐf�X�)���&���!ZQ�z]&�����}ݍ�j��C�tnnf�N�k�����j4='�N� B��&@��?���bbI��F~6=Kԙ�A�p�x�?�9��L�h�E�E�ʑ��̵P$ݏV�bd�Xw�X�ƪ�{x��Ng�i0�Yv�qw�D̤�F{���6���a�t�繌Bi����������\,�X�(�� dV�wI3�Jؼ�5�g��?��B0�V�����@N �� {t/S��>	r� rq5l�/
�LU�[�,[���K��)ۻ�dP���o��l�Â08ޱ���K=:P�L�\N��,�EՏ��� ���w;���\X�^��0_}�¬�~��!��āG���({�6�]�Z��e�J$�͝ڥ�"���#�y��߉_z9?��=�>s��G��W1�}�[FZJ���\}����Sq�����sK��q@�ORO�y�F��1c ��j���S^�~�̄�tZ̈́-��h5F%v��au��	˽�ci���?еa������!Gym��$G�DOQ���h �b�����y�>���Y�h��-�" �mF;<k�>͆�7��莂�Y[����o�k9�E��K#�'��вM�R�ŵ�����3d�*vVASl�X�b�@��9����a����
X�����彏&���@ف�=S�ui��V4��\�t�Y�U4�t��]]�S���jc;UY�l�t�;��=��ώ���Y�
i�;(l�������cP�R���3~�d*@�R��<��^M�"s��!b9_�~j���V�~~w%��y�7��|k���K<�c`e�
�՚�0H�����IRD(��TߑJE4��Smٌ�dY��c��d����U�-��%(BX�(�Yn�]i+q�,�^���,�=����h�}��
��M�c�7�5�Nܤ�4q���.�0
�|�{ɠ3���N{�m�J�ɯ��!�8k2Y^��S}��f����R� �	��u8I9ЀY��F��h�����wøڗ�h���;Z�4������5�&�τ~d�����E���&b�O�,���k�����l�5�n+_�<2�ݝr�8�C�
w*hH�wf��_���{j��I�"�)(��t��:�V@��?��]���Q�H�V0;�I�%' #��ޒv֔��"r6,=�5�d�i~nTVwU�i�:��H�P�H�2����'b��/�EK� �1��,�Gm�c`0���t˘��"Y��ޅxK������[�e���ɠ����ePjy�Մ˒I��ߊZ���z�Y$��%4a���%<��r�q�8Į&��KOq׉��	�3��W ���H��XZ�p�o���ẹ�p!�\x$kFjվOtG����fB/8z�������T�.�r8f���s:�\�O\�]}�̢HΙ������Kh@���	��m��@���P*O�+nHwHY��
Y�m�	@�q�e1���#�yל�?6&�� &����������+��[W�H�g~h�Չ�͝��[�Lr	�k~�I�3Vl�`��{OX&6YP���Ɨ���	��ۜ����Q�/����i�����#�4�x�ܝ��P�c�L�i����D�	����}�U�JV��sZ.p�&���C(3I����u�C1��?W��F����p.}1���o��C��7���y�DǬ������'�kG�h�@�.���n�{6�N��/��uo�x��Ԯ^uE�L��$[����t�
9��@T� �s�5K���F���(���e]ZA�M"�&́M3�E�O���n�r�l�7�hαܩ��_/���W�b�t�S��UW9�`���/ �wU�{q)t]1"5���i0�cִ>3S4�?n�|����:|��ikJ�Ak��N�1�e�:�C��׹���1^{z���	4��1#��^�IB$Ҩ�|����6�Kx���O��Z�JJ���aFV^��#�*���r��EK�f�@`@c�tnn�I��@���J��������t�i�@$��:����#CN�C_��{E���C	�1i<툋E�L]<͍:�~�,�љ�a�G��G�D�4WU�q�~��*u�;)0S�C42	��U�̶�1��5�m�P>�ê Zz<�%��eF��IM�
�r�E@ɴZ��H���z��,?�ĉ+�V>���ޟ^Ɗ�����ۏu�*�W�o�%�gn���C�N;��u�HK�Hj6����:�K���E1�����\~�Т�c{����=������Z�Wo�@���7�����e�"d0�iv�x����.Z�dr���cf�7(+���W���i"�#ɹ�-��r9�Ö�?{T��g���)���%+F!nnm�s9�����1K[Ȣ�5AK
Z ���뚋89WߤҺ�CU�.�W��`�9\��;����Gqv��ڳ�_���L��K��0q��>�i~/+�";��[��`&�#�4ќ�騆���5?,�&����(����b�\u�����f����v�p�I�ڿ9(�M�4P+�s�:�'"�NQ�:��1j��L������Uܷ��e��@Z�l��Q��L��� 3�idJ;�%��"D���1o��I_���MSX6���ۀ�����@�1�q݂�h���Yy��a���κ��c�[_�D�d}�(:���w���z�* %�����U8ߨa��L_���d�hX�)�y�_ܘ��[ٙJ�d	De��̨74����)� O�������Q�U�&Z��?�j2��� ���GG�q�&Mn-��o��X?h<_Vy�'x���5ދ<��N�X�P	�E�n%�2g���k���:>���O��|۾�����[Xq�(�b���f��]�aKi^u�"�`�c��J��@��|\��~�l/0A�}R~�[e?ə�Äg��D$N�[:fB��d�^����'��D�Ve��ư��c-���^����|�nW�p�l�Y
�i.y�	����	h�H2g�<�l�>�:X���n &UZ����r�q�y��Ч��\z���(>/y����O��͢o1�Tz~�C�A�:(��)�*� ?]�^��E��=6Bdd���p�����C�YA+�l��UX������Y��6�?��í*��c��Ǘ.7���L���r�zP%1'1� ���q&V��/�@���9	f�C�8�S(}�w���0ʹ�JXJ��L����m�)"���N
w���	i�(�V�`�z��l|�ZSAs�3��1h^wdd���Rc����J&h�ԑKAT�tX9��b��8��d�C��/�|!T�F��olȔ�m"P���]ǫ�a9�Y�[����B)P��0+py�`�� x��ofƐ{�����/u9�n����/nN~5��3�}��*܁��i�
X#|�����j+R��Mq�+Q�8�`�����A��"�H��l��뭆�7�v3�u����u���v\����\�_��̤q�~��TDD�)�����$�=?y�V�q n���� �bۇ�>��L��Gѩ���~���G0�W���, ���I=�\vQ:��@�xlzxi�>u��v�<Ѕ\����#�ْ��3˺i���uPO##}���:�`%�$��F�e\����{CTb%�����t���-����Ş�dT���_i,��w�-'��l�%�#7�-2��G����h����cUjS�RBs÷K�P��|�.W��� ��#[<q{�!�1�,ʶ�$��N�F� ���E�0^�t���y(��v��X��q�FF00�$a���)�x�d��$WB�B���؁(,�I�.����rX���#��H_���ʁ��p��$4.�*�В��X�>Z7Z>�4[�Vo���E��u��T�W_ą�|�E�\�Kw�?���m�^6K{����j�XTwz��Z���Qc��2������Apa��'=5��kb)ꍍ���Mi������CGm���"u@��Sڭb�`׀dm�
�UJ\͆��F��／� Iy�3>~&����ɚ,^��v���6�/���@�.��p��n�{�B������;q��������sKt����"�sL�4��H�%���ǲt�����/����e��E�ܖ�f���6R��Y�{	`�S�![�r}w�o�aڅ<���!��]����	�D+J6�bYg5Ƕ<*��3���M_xN�}������>'�hf�_4�e��-�)��O)��\|'�`�۾=i�����U2��=V�(��щ��f>e[ը
=����Ʈ1@��VG׮p?��:ȃ�jE9X��ZO0����$r8�e��������iԚ��`��-�� j�vn�5#,�u��P�xSµ���������E[՝$v�O��*��f3�1�U6�(-���]��j*����ď~j�̶�B�p�wX�4��Z�Q)�+�Q��oOV"i���ν����I0��~��¹����=z���g���ph넋���n���4Iz��W��k�����dT��!����� ��e'��W�px������x�����1`"m`ƪ��C�Ƽr�x�$�b��%�EH�>r�����9�0���xѝ�z!�:�zE#KLD1~���2��J6	���c�ŹrĬQ��w��b��z��*4q���z�����VF��9OL�rI��v�y�2BޢVt�`.]fQ.bu(%5%�{�N�.� c������u�(��]���dwc�ߣ�(;�z$駏7ұO;���/,)�/�'k�A(��Us")�IN����x`��<yWX�^�[�&�- �㬪L���_+�m�_����0�z��_�y���K��=���g��U6�?C��w���A
Ww����2����%�-8hvlc#�EDw�{T��s��6ة`2R��H6����$�C�Z��u/�Uw�F��f�@��e�����/��S��g4v����{�ߎ������kjJ��O�|�R�3�8C��Q��WoUg��7|]�̄3@��A�=��5����&5x��QXb�� �]TC���&~IO���TKmKZ5��ȣ��xz�r	�}?,�T�cJ�'6�~+0��
��� �l��ù��������3;7aa%?�TO���	qE�Z�0/�۽b@�9}������v� ���JC�V	�>+�y��U׉���0]P�ϯ���+%��>_ ~��$(%Ӝ�*j�����R���|�և�G��91��\�4�1�uN�ے�exׅ���HV�πfA���*���[i�G4�!�h܅N���n�)=~�X�BWj{h���}8W�M�c�7Zb���T_���lp��x���������/�E���EfX���O���0�MvFn���*�!t��,1���5�ʐ��N�5W�)��D�O8��+�!L���n���cL����ow�p� ��#�?Hg��by;6BE��xy�h}���CQ��33�e�ͼE��Ы��� ����a������s~��(�#���)�bECW��$��m����6�˸����5�j8�d��)G1�=���ޥ�\����D�N���P�(Y�S���mn���E��J�pc{�� �\�Fp��y}�b��P$�CeZ?.�I�����`X�1��R��($�j��u.�`䎃ȇ���:�Nѽ����mg�3�ԆC�:�����w]î�p���7���Ă���6IǏ��C"���������{���ln�`a��Iu�^�{��@�"T�t�x�t�\~`�Y�| ��D� ��C9qF�o[Ws�D���|q�M~����ʰ���I�v��l媣�$�s��٬��L}�������g��+8K����w�!̛�\�%���h�&�W�\���!
��9:�/���t*�$��~�k�l`_l����q�~�l�e��7�ra}�6&A��7����K�
�A߼�t�oy�D�+r�T����r�fS막e6I��b�}��!��.��_����[@�x@yLhJH�4x.�Q��dSt�<����D�J�a_��9y��aGy$�^@� �sK�Q'���t%U�t�����_L�pȍ�P�cs��Z@����5c5����FF��PH��O������K+�bQ-r�0⬜�I��{���[��)����@�PYP�\勇�b�zn8�&j�;	Z���X��M��ص��Q��d�^	�^10�`k�fj����P����hLb^覙
R�i��@���y#�E��ٵ�\!"ǉ�'���=��Fd[��IД�֎г�[�%H6�ҖQ4��I���떫��g���'�ؘ}���9Q|����a׉�C�?���h�3�&��Vst�$b��C��v��ܲ��<���
@NxPP�"�5���؉�2:�#��ׁj^���!f��@�����lh�����6�RVΝ��L�����T�6�h�8]6/(���#i�A�ҋ��N� a���g���£�@�Ӵ!')؅����TTQJ�>�?�s���`�4�����y��L�T�*�Ӎ��
:��[�9���"����d~SG�fg[Mb�U!����B9>G��x�jZ�p�q�:Z�HL�V�v�DPף
/��;ߢ��>�R� ��v�����a� o�7zD�V�ާ�x����S%�V(�+O���<'T�8�L20f��Im��]LSH�T������;�FG�A�,��X}�,̈́"u����HM_�㮽f1�9A����3�.�y�_�Igh��W�li����zq	(bqc�\H/��w"b)@��n�j��fv+l�ـ�q��*VI۴�i<�C���D+8N��Ȋ9z^����t��=L�=bQ��f��nڕ�$����x@U��p�����`]x{����:x5��tڊFS�TA�FB������b�� M ��^�z
j._y�|Fβ1��m�xK��2�6Xs���0pJ����	/��r���^���i
��y?0��}Ś����+h���H�	f3:�����޶��:�dy��zv'�7a�n �>B�' �v�I�r����!���+١x�#z�@pB!&����b-��r��n��q�6����u ��#~�տًkb��j��o8�
�#^mڢ��5{�VZ����J0�T�b��r�	D�sG�G������r ���l���JG$!�M5��� �$�Fi����l��vR�_����z@���S��N���L�8l	��N Y� Z�2�Ⲗ�f3��K�,t�F���J�4O2��[�����<��Ocx)R�e,�vsW3��m��FG8����� _.Z��z�����at�8O�QU�c��nMnA!�Z�n�'�q��m�F���X��?���oԀ~>e��.��N���0��I"S����A��6^5@����&ܳ54�sBtt@3d���0��h��§?e��cR�-n)_�Q;la_Ah�&��Q�
gC�7��,�',����j.eo��G5�'d�P�'943���4LYu��b_����Ґ�������1�C��j���oO��1�I��}�󪣓�!�BQ��!b�[%�2S������*�Z���p��\�R�����g�1L0����s)@6��Iܠ���j��&e0p.M��0��5�I���;k�������Tk��~BYa�(״�֚���W�iq�8̖�"�	-�j�]ZU�Jy�����}���1���g�
��J���
�[��������i;�֍f�&#�J5��	�L���>v�-pyV���o~f3聰�6%���5�:��G`'Vdl&���ҳ�����f��L�Ѕ��"ג{��P���{��e�o��+m���3���P8?�Z�V.*�\��_�巉���ּ���f��C��>��nmt��.5w�n�l5�C�Lp<��8��[�V����\�0@A��8�f�,4�2�u�4q�e�:0G�6e���r�wI��(hc����������$Ϟ^�i#o�YS^��]4����_�e;T�E<���~���xi�Nȍ7���}ZI��@��-��q%H���T:�y��$I���1�V����	VV6Y-�f��:I~؅��E��oVE��Q�7��x5^#�4>`2J��z��E�h�M�l�|P�G��,��;u ��V��*Eƺ�1�P.�mщ�*_����v@�'�h�ŒA����G��t.�ԷX��=�2Y�mWA�I����ã�:`ֵF�C���6��u w�.�a�dI��b$�[ȥ尿���Ͳ�[=�#
�!@��oόf�m�:x!��?�N�C�d s��ħYMI��#�j�|/V�SE{�1�-<�vY_"7^B��SB���"��4*���!��Ee'8b<�9��}�����<:�^�RWgk�Ieu�J�/[��{��dC(-~���I�@8��Qp�����C!�R�SJ�\�
������ԸE𰦦馱�ޔ�� R����kscr����F'nF+H��ƿ�A7�7�yB�Q�u���h_�RԄy<^.g+K`W>�MQ9_G�M�W*���6j Kؘ�W����(T��\z���ݘ�L�6���w�Pq
�F��.�?^���N��5�7;2J�ǏP�`LĂ/Mܡ^�-w##�0�;Ͳ�| ���
w|>B㔮G�j� y�Q�oS3>Ǡ"&]#�Xj/y�R�|��1�k�4�U���@��o��f��R)pl��.��vFa� <U��{��	Eu_rEe�̳����-j�Y��6�:&��SƂ>��Qyc�3����O��r�	;%<�&�?3Y�l��#��~	"��~X�S`�7'0�Cwn�\Rk���1�,��W(U#̠2,/��)Z��g�9Ђ�18�?���D0�1�=֕V,�(�;�[��HGH�5c@u��\��<n?�4-A����a����X����kf1Bg��T��A����z��ۤ;�����$���L�Zܨ��ukYÜp�����������P�L���He��!,�]�]eP�rp>��=��r��{���UeI��؇=g�:��% ,�@}����������߅6a8������$�2<U:1w{�j��j+01	�����I���f�c�y@��v
L�`��W�6�Q�U�16�*�/��I�-�{ɴ���8��'�ms^�%k
��T��0�ܳ��KJ��KX��n��	 �Adc��e8�#OϦ��jal$)���^����_����[t��Jz��8``7:t�I��u�楇��W����9	�yN�����;���Ҏ��'Cϲa>S�)E4�o�1<S��!	k1@�v��E2&I�?�ePg ��A��*�7��-+�%���.�<���c�s���9#�9_ok�z&��W/Qre@�r���R'��^��k�ZV�I����K3���=K�ϑ���R���K�}��41b2L�5et�+2���&ĥ�zM`U�c�*oF��� �"����<b�?B�.�"�زXk|B��i>{,���¨������%�4|q?6�_#��k.�e���Vg��2#�b[(o5�
��jEh����V�ݓ[l�'�[���)o�����,��m�)�X������~B�BJ���t��Hala����"6�!D����Au�eq�x)�Ӱ˧�;�׎�b�.5��ֆ8Ɂ��ã��f�@le>�zc�?:�PC�0��_��vE��5�B^��]OE�U�`�WLըC^�(�%z �R���
_$���ʙ�B�ٲ����q���&� ���
l�R��"<;��O��5틣Y_,`&��d�Y����g�jq�Pd#8sǶ�VPYQ�C�	�C�۹ Xr(hf���+�#g:v�C����UP��s瘁X��Z���<�oa]��ШocO�����nȺp�{��qy��DٙP����]���N�@�pr,s��zb�0�a ��iiWٮ��n=�c�⳪�5���8��S��y���*&#ohv�Z�����?�F�<�������2V�9���E׋��n"^z�M�^��e\acSt�s,"�L�S{�mA�9�uQ�1C�hW9M���f?�V�a�Nj�h/���C����GG7��O<��*���,CHk0��M�i1��'K���#���:1LŽ�ֈ�E4�<H`�N#��j�:�u�7������æ�w7�|(�n`+��������R�F�Z����n��]�\C�0a�������џ�C��q�(�rY��1���c�tv�t��.�^"з[`�g�p-�@uV�H�%/���� Z��'����14,T0C��t�eR���Q���ſ�Rעh�*��E�U鎾@ŎU%G*"a�� ���B�r�{���cj<z��Ae1fe̯�3����̐Y���/M<�ȣ��#k��*�6=���h�[�|?��^��,rd���VZy^�g�qP��O��/!n>����ȅ�'�S΀���rL�.O�;�û<=�Ħ��
����PL��v��BlCU%��	h�>��W�#�|Z�kW!\i�@�s�3��4�W�$BO7s�H�	´�t�%Q�}��'�%����9/ݐw�GN#�y�q�$����u"@~sh��XO�?o��4bP�9,L歺��ƹb�j��=��r��&��������)��`^#[�7Y�Ab]O�uԺ}���tWl#O��+��.�'=
�B�A5~�Yc]#�7�vKF/ʯ)���J�nJ~n V-�1���i�8�XVT��2l?��MΪ��xq.�����1k��Np%��xC��7�ǝ�F�&K�A�P��c�û�h�5�o�7�lt~$CH�R�(���=D]��<o�dq�<���*Bp�i��f��=+kϚ��Yi���AB�-14��F���V^��R���L��m��[OQ��$�g狳=ѫ�hv�W�<��)�>F���Y6�	UN����:,����7Ԓ���o���"�6�Ỻ@x�Cm�����Q�f�/��!ә�$�2�w �$T�8n�3^ɚ�vxTr�1��k]��I�YvZ���[\ʕސB/�xR�8�'M-��P��Q$� i��`��q�U�suVy|"vMl!�%�?3�Q*A�-�5(���Ln�N�8"}�]M�8�Df=�{;��.f�@!�B���[%���9#����j�C\g��W\L/����L��3�A�_�-�����/ LI*ND��1����7��� r�Ɔ�ŊN�>�.���ө���/��r������q��t�o�L��6�^g��,�} �<Ļ��a!��^��'cZ�{�rzX|�0�*q���8������yL�u�Rx~E:I�G�u�)zqevɠ NI�SQ��I�����8����,����i�����E���քbdW����+�ڢ���H4rհ��y�^˓g*���y��m�\����U�l��gэ~l���}�������(���c�}ͫ�1M���N��n|c�M���n�[�����[S��@)aͩ���������%z|qJO��ET�.So���TU)C��n�e1���5A�m���+d�Z�O��;$Ӷ���a�n�S�e�Kz�3�H���$
7���n�q&"�
���wh(����+�����m+௧9�V_�;�y��H[Gd��-���� �*�-p7ֿUr
+��/N؎~c]$plKJ��tQ���k����+r���V���ΊyIa,t��D�0��C�����E����:T���й%�ep:a����!��p��E�e�������i;rJ����l��-�ލ����f>�M�@�=�%ş?*�+\,��tf�a%D椼�|Gc��9*��RM�A��t���6�`ţ���.Z���ּ�/1 YZ���F!w�\��TI]:r�k+6r˻W���\�ߖ:�b����$H��	�svƵ烑��6���vdX�zEw�7O�`x�L��[uX!��q�\�f��iś�|��],�W�>M������'��,��VK0�R�9�#����=���G�굵,Y>�\L�T$�n�d� 07�����n�dH�]�c8����&���}��)�Wà�[#7����x�O4ZkHP�LŁ�.o��f�AA�8�\�W�����Ւ,&�<2���h*H�D#s��TY$o,�L��ȇ"p#�A�U�t��{����b;�;��:�+�U1Ԋ�W� ͙NT��{�gθ9��`xJt9 �s�2��>Q�cA�ҙz&�����1��e>L�$�{�|�E�?0��巙���~)B�_�%>������_�ԣ*Ät���[7���wB�,Ar��(���4�wڒ*8���;T�0�viw ��N5������)p?{�u��^��2XE ��nދ�bھ�������Vaͤ�B�O^rm���̧�����@b+[��I���	't�Ƽ@���vj[h����U�2�AU z7ZY��c��t�ǌ�C=�n����3|���Q�87.�g���6��}�J~����y�4L �FR�iЅ���E�Q�CQ�y)�3�km��V(�rGK�o�{��7nj�Y�lAw:��٫�2�o�B��{�
;�֮��~������
q�m���/yn�q��cmi!���W���)$����ٿ$�I�B��u�0��x	2�: l��UvkD7����V�vC�1kb���]���(�jM6�撢�1T�M8C%ƃMFF'�~��nQ��y'�t���#8;m	���|%���S�����.�@Ѳ�]A�� �Gk3<<�63���%=�h���֙�4������4R��`"4�ă�W��W��2�ꬸ�I���0� �!�/,TY'�R;�Me3���r�dǅ��S\�Ȯ�%}�hf��@��8��V+���ҸWesR� ��P�+��m�M��S��'.�aƐk���2i�w1��rqz�9p^IU��v)��yW1L��`��B&&�_���7�x2��m
s���Axa�q�;�"����!i�eeal<�WCDZLΕ�������u�ߖa��eoa�Yz��s�f�yP�B3�~�S΁@�ɺ��1��s�y�b�NԾ>�<��IH������{"�B���=����RYG"f�Is������pH.��w���ӏ��B��i��}Ob���w%��\,*�e��K��Ɍ�K����r�j `)��Qt����K��8����lsYVȔ���Oʹ{�f	�b��+�����e�=Z�$�4KS�_?b/��4Q��?��f�}��au����Cօ�HL�W@�TF��".H�}/6A%~"B��V<���~�K�yk!�����x?/DqA;q��JOQ��F��jP�۽yH�'ȫ�W��*���*��,ۍ�ZG��_�m��B{� �赓�7�5؏�V��Zn_�L�̅�MB�7�F��iͯ{��=ezk��1/�F�����9�k)u��B0�0�s�T��´gQ�>q�t�����GY�ZI���g"k"����@�b|��ҹ�2��w�E~��@�'w&`���U���)�:�>_LU�:�)�'�v�����S���m;/x>F�eB=� ���^����偨Y�DD�Yi�Q���ODs��>;����$h��5i�X���������Md(B�j3�8��%����cW�;_��.�c����1q����>6���f��/�"�}��.���;h|��Gy�9���S���Y|�+n�m��6!��O�sF��W�fh��U�g}�-=h�@�}��Z��H۽�V8�+�6ڗ�w8�$;e���8�����OߙBs�g;[qpQJJ%76&^J���f�G��녧�B\[mnü�)�Ū�6���B:���c$u�i�v���~�#�@�Āw�~����|}�����E2�XzX@��g,�ŷ�*n�qͬ��ᯆ|CVSm���D�W+�r�٩��f�SO��s�H6A�W�c��Q�}�5��k�i=S��$U��9�l���D�)c��+|�w�#*O;�T���c��L�9���_8.q9���_Q�J��󦷕��p�u+���M.����i�Q�x6d�&��?}_�3�%���������Nhy��{�=5�LJ-M��>��JL@	��yG\8�M���#�������Ւ��t���!�vh�"���̄|XǏQ���6�Z��	X y]���L��{X��V��eT5���r�g-��̻�v}ߠ{�_�Eh-{֌��S�.JUv�fMv�����U�)*��As�T޳��<>��]JG���W�*YD<���;^�+j�ώ!�iQ�����(F	�m�g��}��O�h�Z[Z�Z�?j���-2՟j���
���ȯ2F
!�p�飧�=hʌ�E�C\�4j���*^R/�wZŪX�I�B�2V\!�#�+FF4�?��G�	���� p�L�%���&�,$��?a�џ`p�[ �+P '���%o�x�l>�\[Y�%8�8����!bqڊ�{����B�=~f<��Z����u,�d�I�3��veqm�*�ش�r|,*�ܷ^��:�f��Պ0���}���}D�W�H��j;�K~�>��_���M��jt�x�t.�3����l�y� �z1]t���v�.���L�v]���xn�:>�#��"�͸���ex�AT�Ϲ%(�K�"��t���d:��.JUs�� �Nhr�O��C͍�ԐjQ��NB�?�%=o�6lH��������)Q~~�y��շ��g-27�*��h������N$���S
S>nb'w&��+L˛��3	(�7��a^YTS�R�$.�n��ѝ��N��u�3��Jy�r���5�9�`+������$g��� ���=���=�c%-�I]�wd2ӄ"�Rp�ɂ��P��(^H1�8��Y��C �1��M�b��G��(q�t��!��w�_��iz��cн��[O�h�9�D~9��1��(V�ä� D_�i����iG��>Ŵ=�Ih[��o;���Zpgq`ӗ�A�/c0���꒽� ���(�멿�#�}~;'2�� ����9�]��v�-���Q�
U��h۠��9��b��)��^my̰��)�r��.�<��q�[ Æ��Na�{]l���ò���9U�Al7,�ތ
�sz���2�)��Jo��|�%�"˥��O�r�K�H
��yV� ����G_A\���鸇�g&�U���\.y�/a�p��Jt�Qd)�W�.�ݼ{|a�o������˰�Ɔ���oE���0\���������G`��<�s�]��50��V�č� �;i��˚z�h�Y:r'�3��%�v�p2E�
K�����n2��"]b��C_���{�e�������F�|k��7F�N�J0T�ܾ�t�}hEQ��5[��r�W��GIc`�d��	O>���7D���/�ZA��Y6�<�� ��8����G���l�����^������G|��)�L������HÄ�D����ubs�A�U�g�ҥ��\�h�����l��V�oTD���rK<9l���%U0�{��G�gM�by�QS��EJN�R��]�?6xpA!<�� ���͏��Hi9�>s��e��vR��g����!�Z^E��?�����H�ntҤ2��{z�:���� (���3D�@�bu���h��/mG�(b��wj��î�ͣ0�R�ﷇ�_)��)�'�m�߉��o.�:p���k)@����K��֋�es�8����dty]Nm�iG4nԘZ�ha��1��h&�yxv�����qҦ�;P�P�A�����ЕJ!\$�O8��z~3���n'��b�G���'���)�.d󌲙O���9�[׺��Y\�aQ��c��\�@(�^/��X�����	�h=�Է�򖕈�u\�w����$�U��KC��^��������H�5oI^|�Gű��=��!��QZ3�x^���w����.��}��o^3SčyW�T��1uX~�/�ړ�C ��K��t>e��K���i�`|�UǙ�kH��̩K$@4T�ױǨ��!Uw䶀o�)\��vUҬ<azrewJ���Q�c�[�덋����3�oS8\b��q��N��W]���9J���1� A�녂7�й��$孽~l���P�0-J�W@�`b���ZR���	p��AD�K���������`l�;�����ἳJίG�C��3}u`��i��@Wl+	�='B�7�E0<��S;dmy�>����'�>�\����s�~���B:~q�����Ⱦ� x}�ek+U�%5��x�7�<h 妸#����F�7���a[ѓ�M_�L;N�0g*0�SȈ��鬈�:����z<���>s�o�Cx֢�����/�`\�Y��۲���;3��R��n���o=Q;�{`tۜ\��:ȳ�����n���SR�Q#��նs��q�-��x��i����)85���5�ܟ���*L��[~���I����ҪF�ԨE 
��_�~�|��o�Hi	��Y��W�B���K��Jc���Tg=�ڷ�����FN��=��$JrV���R�@��t����Y��~!�NC���c���ܨ��*��GacH��*ʧ:|v��&s�fE�%��bL)Y�j��3{��/����P�&���$�6��pGZ8uM���PS�"`�s���Z!J����/�^�]�����?2^ڸ׻X��~��Ϩ
�k��$+]�tō�y�jxG^%<���b�s1���@^?���S=(�D�h�3���UyH�̎���"R�=s]ql�̻ưA,j�_��� q*�+Ȗέ��e�����JV%�9{����S��yE�﬎�?6ezRC �[����p��0bV�)��fw͘gO�o(��� �,	Zc�v@Kȑ1��>w�MiXǗ�LB��O��iG%�Gd.HK�#��Y&��N[Q`MZ�i#p���|����ĉy ��� mI�j�E�r�<w9=�L���$��7�@� ����j���s�/`S��3����T���{[�W���K���3�G������C��#���QŔ$@��)����S,%�b_nlD�K�J�g�����Ď����7��Ѧ̟5��wZM��/��Up�����K�X�Y���&y�����9s�a��*1Cٲ��O��־H<�q�OsJϺ��v{��E�1�tɂ-�����N�{�OQ:�4���	$��o~Ie�`mU�_&2�Z�cz{���"�5TI0���rG�GB��H�F��]5�1qE"ڲ`U�҈�,��??��-�/F#��h��Ό4��r�J�����Gu���m�.����-*=��+U��T}"�
��ʹ��;�����#v`����&������NLZ�em��M1X�q�:�d*2��&@I����EʀI�C�a�za��h]؇!�AF��zo�rL�{�@k�lk>W��]P\O��1(�b�����^��eSa9u��,V��Ǭg":p>��b�72�Q�l3Kns�>���G��g�R�n����*��2?Tb�J)]��*��n=�#J���Ѧ��m�_��&�58�]@|飥��3uY�D�"����948͂�aB�ex�"+峓�}� h�����ϙ���x(�<��,�����0��u�;��B����P�HZ#؉���M
�lH)!��}���d �H#_�D���v(m�BLe��#���R���_�� k�	$.�mb�nQ���d��qV1�"�~����M�{�VȌӘE{
]o�bl��:�k�	��|e �M��0%�؇��d����ހ��Yy,����{���7غ�P�`��Q�� i4G|&��݅�E�3�n(G#W��ϽlYH��q�Ok�1>�ZQ�踫���2�+�s��p"�>&�xMR9"^���o�D��(�T�����Komg�h&6�{����7���T�zf߭y���}C��W�~��p��m4�a$0(���RB�(�{� OhB�8ͨ�X���w�0���[���J���K�>����U�r?���
�$�ڄ��p�!7��F���ۘ����Fa��'��,$���Y8?��E��qh��j[a/ҡ��]��+��r���[�I�\!�/���E�YGR RƄ���SF�.f�n�~ɮ���s#�Y��RA\T|�OڏM��nZ��~e22()�̛�w�EO{���P��/Z�l
e�&�T+��3܋ւ���&�6�&�^�*�a-�v�:���ղx(��#����o��B�o)�X�,����2����<��*�g{��� ��2uЭ$�7�O�K�zW�ُ�$��mӟ�� ��ddӛI�����5G�P��xbN�د��C�lm��G)�-���<�e�P?�I�|��:��c��L�䥚>b0�ɼyc"R���A��p���L�flw�঳0��ʙ�)Ã�"���괋��ws�b��J��I���i�87�G���&�N :�ܖm�ٌ���-k��MU{��)�d7�|kݥ��=X���}x�mƆ�D��=J ��z+Pa�c䜇��@O��g�Ü��.��Oai۳�\܇t�����.W�.��
s%�X���0�|Ќ�����[M�I�p)uDU*j0��|Uv�և\��J[R-�gp���&Q��f�^QRg�=��9G�h:�of��҆5~]a��lL8�0At��(�݇9����p�W&�TI���J�o�\o)	�'5 ��/����I��X��>�#�
UN��G�YG��(���xi�Xz�(1הms��/J.�-x\3�]��bC���jfq�/�Ox�����l1�z������y�n�>�ʐ��٨�qH^q�;L욡����E��H���kr�0brӲ���]1
�ӈC.{��m���I��̭
��ö%�R�f�B��s��D�ö����ϰ��s�;h���۬ޤ�'���.w�Dr�3yҩ+���c![�P�P[}5��D^�"$1� N�N�V�cO�c��`YHó�z�?r��y�+9��Vh29=����kBm��G(G��)�J�p#|�|�it�1�*�kdcYE�����:��0LK"��t�¬��ة_!�ڽ�:�-���H"�Vu��}����L�"�����ʨ��Y��|q��{�FFo<�q�s��v��+u�
L�}[�)Cf�U�����*�m6�%�R��:��m̭������[�D�z"c�@{\V�vIY%Ԕ}Fn�L�`�p����a�Ƴ#9'LS�@�;�=���d2ҏP1�eeH�a����?s*¦_�aiH�z&r{�HQ>(-�5�d�'eNHylô�G?���z�=C�4X}J��c-4��s`��x���CB������v���S��,�]���c�,�)�4ɉ�.8<H"�W��Dx؊5����U�O��;t}�����yf�F]d�'��P�V�=~����	N��6�x7K�.�B�Ur;	ou����:�⪌.�(݃��wЕ��w��j1(Υ�M�oL ���oL(+&Z��3�9��\�%�*6g�'Ԟ{-+oDA�❨����z�&-5�-Q����ZNQk%d��YJ���@^�3 3}Ŕ҈�L���bz�]fWt� }��a�Pܮ���b���Z[�z
S�]����\@��?��{n���%@���.{�vleu0@������R�1Zl�[�C�ц	Ւ�h��{��ϑ�ɛ��RdZu8*X��x8ΟgQ�ԉ%��>�1�?S���T*{���T'*%�Pbܧs�������f�CS)(@ j���mA��PEpT"��� ��u�{YA�c~Fʵe�L�����y��5�(�	�z/"z���*��6�_/9nu�H3H����Lh�'�N���e�?.w��@-<�l�67�3��|�=���$i_��3f� 9�o� x���1�h.ƴ�9V�s���9!Ȋ��ȦF�A�]�7�,�߯:Z�p<f��3ĥ�˿�aHbxQ}��k�wJ�á��f�*P�n�21<gi��j����.J�3� �Mx��~ :"8�������a�ŏ"�J�/�S�? 
�c�w���9�e�PF ͣ}�'���ouc�g=�@�x��3)A1��I�{R�Ǒ��[;�u�-���6%c�.C@�οK_gv-ߌ��Å�V��;ms��h[=�?0�0Q��y���q@V��M$�Н�S�2�N>Z0|�3\���*>���(D��D�4̯`�ɨ�˓�*���O)˞o�D60Ŕ�W��l�Tz������1��ʖ��i���x�����1��L ^_-�@�9A���R�W.�"C�v �N#���8W-=�V�jf��?����v͖�׫dGٱ���^��3�9t�J4(���O�aIv�^�m�C�f!�p��������*�ت����E�[)����g-~��7ܾ�!26I�e^���� .XI]0[w��E�p��[3��H1\`��Ek��¨��7��v�\��f�2���鹡��Zv�D�$�(��K3��e�s!3*ZO�E��/6�2���?+��z��1[��ݘ�z35�-8F���s�!F����̛��I�C�)���P�Oa���Y���|���p%��[�j{���李�?�A�~!��K��x�ԉ��Iye��`�r�:��T�g1�gA�%��s�&�t�ý����'N�'�W���_,��X��MP�+�$��Dft�{��;~؍�5f7�us1Eh�-��~Za=�s�� Eo�N�ܫ�R�O��ѻ{H�9S}���wk Doo�o"����Dy�����<o�4��� ��@�u�P?�Z����i�g-s%5^\;��P� �&��%x�N��2������
��u�Ό@q�ׯ�d�d�������nll�v�����s��6C�(��jvtX�W�2Y��/�lA���b��})z|��)y��Y��K�ȹ)$�%�p rd���M����H�0f��B�fv�Z!�@�_y�Y�֭�%��P�/˕�^���ә�����d���֒V���^��7d⦜�#�beԄ�����ԋ�����o�t[[u�g"l���m�$R	F�~U�3d�C [z����{�rI��ww{�vV�A�}��t�C����9D�Ղ�ڠ���<��������
��+{�2��/��]D,�y� �ZnZ�Lz6x�!X8���k�J��I��q?3�H�<���Ξ�ަ����*01Poܥ�����oˁQU�J����ka�otW�U�^�������d!,����$[��H6��AEc�,�O���N�/o?m���.c-W{�_=(D�& ���I7v�X�]�PS���$&Ï�
�>��ps�jzaH�<��˹�(8i∅.�t
�B����9BP$���#n�����wVO�T3v�I�ֽ�,*]D88��j�T�?]r�|���FH| + ��?h���0r���O+���`FٿU娦��k�̪´+���2
V��\ኇv����G�3�ec��;q�s~��Jc�<��W��*k|�9?�RV����WzD���A��n]^=�r�Q�ˮ)����c���&	�G��@�#�Y�N3����50�T0Em���Y&_�ۙ4-90ʦȸ���m3��/x�qߣ��5���i.����s;��b5�6�4ڣ����#.��h\>5����a���+(��N��T�ɹ��F��'�e��L�H_�23R4�Ϊ'�F����P+�?`%�ryBj5�Rj�̚���5�a��B9��9������޳$[�^�N�;�e	�_�Ű���g��)6?W]>�(��� ;_��3�`6|�2J��#�4ը,*�ڑj�~]�"�:����H'�5�xzb(���	�m
���{��	��G��r�{iZd0*�w6eHv�	��4�R�a\!���Heʽr�べ�w}�H��*q�5��.Q��bĜ���[���k��z3��bl˰�,�,��\ڬ�����`>�E�V��Uu�L��n�����l�۴��9��eM�q #�T�x�v���[�{/e��a-�G)�5�U���r�RH�#��~�QXuظ#0]fy*�7Ci3�X�ə$�?	;��@=Gp2)mւ�]�@�����E��)A:����AN�P�<�l�z>��qFRu������+���z��p=v:m�V�Y�|%N|��:��M:���.���R5Ѻ���@2w&���ƿ55�оb�y�i'Uw6�Z�BD�͍�3.d�-���F�8fqa닽��ӌ�e��Ul,b�i���@W4���+ּZx�@sF�����5_U�^��=��2f�=\��I-��L�J�@�����{�X��T�QǍ0� ��k�����m�O� �Z�o��@�\��Em��6�3�}��n�bYpZ`�P����ר`i��hjT�f���_iO`��8����{R#� �,(�쁿VXd�.�����|��h�5�bwH�$h��,�ʦ}��?������m����TW*�0�ٽ���M����<��S8�xH���]#n<(u��5 ���xyגO��t����~x��g�cս+���ݰb-k�[�h�\~��8�K�dF����b쫑�(�u��k��=
H����!��� ��e�U%4��*�o!����4O/R)D�cvuM>���!���x�����woMZ��R��\5sY4j�i���R�-:�+����Y��j�V��]+CǤ�<HF)n05%i�&�~�G�elɓr�%�)d{�#{�ytU%�^0��f�ۗ{3	�ӐJ=�e*W֭����|u���s-*O�c��w2�f���cpP��2�&M;X���l�S\��dߜs�i�A����r�{���-���id���8�C��/57t�����䴊]HR$�+��	e�<D�̴D��6�TcM�����eU��Y�'m-�����ET�v��H��D;���qi�pp�~��~�>�Z�#u$C�JD	&0��g&���h9ŬX�-:!�_�r�ќSm��ռ�0
r�*06b���6�C���>@�bo���0�V%����hiB����È��&s q�J���(�c�f�VV;�n�}�Z�Ƣg�����"�qx��%Loudl��f5����(,����!��"���	��c�t��}C�DAˁ� �,���KJ�V"��J�ۧ'e�[*�LT��-����E�|�z��TT �]mW<yg�"�)�W��M�l�9���m0rn2�P&O��u��.<�QIY$sq*klD�-j�,ߜ�q����X�;�"�(����\j���V��V�5�J�jC�����PG+����eᥘ���cQ������z$~U�p��*텎;��������Kf�q�H���.�Bk8���� �PO
`-6�/����{���<�c ^���$0Ԯ�0��*�4�5��<��8����!�1q���z�� ��n8[�HR�1�h��/�k�X�U~��w$��@��: a��&�V���!������F( H�Gҽ��M%����~5#��{F��a)�W(�FSz��,r;~�v�*�}�_x�֓�;�o�u���B������� �&bt�^���mϘ� h'n�!��B`���3��
Q����q�p��zZ	�"�$�d9���	��I��GZ�;��A"15DT�F�lCbb��6u��ħ��Ns�s��ُ�s�(����ᬵs�ȭ�,=�ӧǀݕ畗�.�����Y^��z9��aC��P,�Dr"��.(͋�D�}o�>�/ʨ
;61��p)��ɾ�!�Z�GK��
48�X�X?L4�򺺳���F��#K�Q�,�]3�>��1Y=`�@��cP���G��O�3;Q5\�r�M�@Fg���&�㔪�{���ת�#�-O8�;/�N �uj��h���;'W��s({:���b�ejY�}H�
g%�*��:��粛�Nj�i&󺣆Y����w��X���N�uf��YCC�VXR�?��g\wG�%U�Q`�Ќ���nꝉ�rx���(Ӛ�wM�LG��e/|9<���(������<���Nds�\_�Z�]���Q��Fsu���Ο_��|8�4���*O��*HR����ծ��z������	C����Ùg"U���Y��Ga�;��B_��s��B�MZ�x�Ns�=�w��%<�hD�7!?+���Q1i c�O��->����/D9�`���iE8���$,MmN�d\a��_���ᦡT�q�!��˖�<s��]������a��b&'1o�Ѓ�3 :1~W�<�>7ښ�Jܚ�՞�b�>z��I�^\h=�w�	<r�����g�&CF��A�O��.��h���lJ� g���YV6o�g���]�օ���fQ���m�p}|�ؖ
7�R4�>q��*p�i�K���M�����0�7U�BS�xZ_��6����x�arcO{j�
ꂠ����=	���y �>�~sE������چΡ͸��Q�8��@�B��d)WJl�X0��@u[^�P?Ԙ��.k,R�P�4��0��qS�}eS}�47_�l�[�?�ͩ���LE�����i����p������7����ʉ��.�E���s���˷��� �6ɤ8[���w���ԟ+��>櫯%�����d���x�N"�7/�}\�y�I������m��z���27�)m�D~�0�T��i���͜&I.��6��e���p�>E�"~4����R���3,�a��b�1dD�若���I�G,�i�i���}����O���\��Ff��9��T�xp�����C��C�P�O�]G�I�q��i���X�d=���5�7	J;��Q�jpOT���nn���,�TvL^��!5K<vTίԪ�L����)��q�6õo`��R_�~b�}��,��3ܵ��Ym$k?Q�㎋u,�;��@���8�1r�_d�x��{"^��|R_vNK(�?�_	�5����WW��hC}���t1d{��?��U��f�����$U�^�ixMp�~��� &'0��N��	FJ<����}���l��o�Q�]�����L9e&��ݙk'=�6����Da�lX	��\�9��fLx��\蘒U�$�A���3{��1�&QC4�
R�1!*������1��<���œc��|��n������fD�u]n�3�A�<��z� `��V�$�����u3>"�Ua�cvP��P���l�P�K�8�����e���7	/���#K��Ty�u��Cl��.G+7`�ہV6B���o�����.+X�|z�d�����9��f�M��J	U�4m-��&�
)42� �S�������rw�����f�u����ڎU�Om�?Zm�ON�9�=�[w��|��4PӮqDT��%@���q���	m9��|LC�ӓ,l��?Uy*Ec��<��KJ���Փ�A��(���f��(^]�Xy;�=��M)�_�u�
,h5/��'�ri�����&��!}���:�������bп�a�'���6�'��f�=��E#*
�;�+��^F�<Sxn�#�96Ջ�/��-�>aq���� d��G1���:��j������Fq;�T:l9ǬD�=�g��9�x�+aژ�2q}7f��N]�c�X�*H�Pg
(Υ��%\�[�W\��ro*������hn� ��b6{�͎a��9���p�nj����D����d�5�(�5Y@ ����ي��Xvƽ�q��
�'��R�O���|w�h��3�1_�������JH��^�K;ee/�	��X��í��1��c<��䇍~�o�&�lY-�]�l��3l2Z� nJ?�5�V�UYKbi?O�����uDF|�hh�������pbIe��@2��T�&R�pr��3�˗��	�U��X�3�1��]8�
�&Ǌ�H��+_��*ɺ����-5e�@W���[��í����lex�K�^k�Q �#���u�����jz>�����>i�^��E��Q��!���d�����5���<��.jf����-�q�"�Me(Mx|��`�0 ��c������-p|Q�ou{2���+��%�ܠ�.�g�KŲt�Na�oV�I�����+�X%��Y�'�XN�Ԫ�͸MS�0 CeT���TE�®�X�Iw:��.�	Sk�P�⾃���l/�R�hR�U ����՝3HCe֓�*׬4��yq�W�v�5j��BWi;w����X�ì˿T�S��W�9�W�����i�!Y��DM�>뢵[�)�	<w�zj�d�fK3,���FZ��3��Dک(��D�4Έ隬"&� ���j>�����Y���`r���'�ճ�:Ɗ�^9'�UVr���0BNL)0&��;%��.�((RR�ݙqd}�W��B����9���=�#���'�H�`�����B 8��[�#��#�S;e����X��9��/j-Q�pO>k}/�(n�-��ם�q-�����-%ne�p���88;���~���2����P�"����vI�5���z��D',��jGp:c�`�B��|��I�Հd.�����]����7��r�8e,Җ"IL K
��F���ϰ-����
�"<����'�@����ـ��[(#�+%I��A�pVSG{���NDY2�TPϱ[f��N��5Q�5f����[S���Z��[&�"��d�u�-��XԵ4޳Y�ĢJ��f��/���s���Tb9){B�P��1=�����^+��֬. +i�"a���/�|:�z�gY/�	��e��ƌƵʮ��p 0��p5,mF�.�$u#j����T.,���S��t�I֗І�[8�?`�ٟ#�7Wqs0��re//�ױ#���t%^]c�Ğ�a_sI�I��t�
�	���E^/&M�)�fiɠ���:@:ih�e9>�[6�5�%�]
?,��IǢ N�W����US���1���t���.'|cF�d��^T��~����򈿙鑵`�Ə��u�`����l�$M�&�6�XPʫ��b���c�qPƏ�A��'�����(��6�0�H�ɏ�4�YD��u�ȣ��^p��_����T}脕#XE�ݙ���]���{��+ҟ�&��p��u ��䕸�s�ԟ�3��X�׀&�?��t�g��#h>�P/M}�7�0@iI�g��}DC����|ȕ����[�hf��L����>�/� @(Az�BZ{���p��|����ϲǨW$�6@w�D�/`[+�	SR�`�]�~��;�ㄥJ �.�Ͳ	�����'*�U�v�Z�$���mL}����/�ρe�
�z�p_�1g�#�Q���L��"8o�ʈ%|}��{�`��Z���?�>J�Jpؑo���7�1DhD����}�m�S��Y1�Q��?�c �ĝ���](z�S�M<�����%�Me艕�Q�a�~C��@�y�s��!�/�MGv���ccO$�YD��de�:��m�N�y&�ѢB����__�Z���Z�·Q�H���=��-+�;&�z*�f[���!Xm�b�����1u��@/����S���'����o�1�Q��;8�@�5�5?�Oq<u!!��OJ���&������,��G��d �s�VT�>�\a_|q�q�η�*�#g(��h)��ÐP��Q����ל���`�����pQ��{�`�F礷1V��ǻ��� 3�+��Ru���֓"�����kN��h��	yh|�K��|]���S��3R�-&pP������q>2;9�=e@��3���/��(誴B�#)��n���1�����i_���QE��*py���:0�	_Y�7+ǚ��}��^t��T�i7��6���ЬO������z��#@\x$I_/�@��ea~�w�}I����M�Y��7��,ja�i�]�3!�3M�,�z�w1��&��;o��s�	U�Ҵ�����=����=.Q���<|y����գ'�w�O�8]Pl�G'�{����]�X�ޣ5��8��,�ʹn����9�5��n�&	W6��܋����q�����=ݚ����ѿgJ	�uJJRM�9�Poŭ��J�F:<�\����|�D?�P�Q���y .'p1T�e�$-F{C�ڧ%.`�;~��.�s�E'¬�݌Υ��gWLW�]:`�p�a^��hg�p�bI���-��t���7~�X�2�����A�mz�ֺƛR��B���̃���R3�͢�fS�U<�(&��H�`�MX'n���k7�cY�"7IJh�Ҕ�X�T5��]�iܱ�Ǭ]H�����-VJ���Am3��w�ن�
�i.8�R��@Qy�Mk��so��3LԴ��$U���?���W��@�4nB�Cm���]
j�����z{��c�z��td�c�Sz�6L�$#������-/���l]*�ɐk]}�	�A�ƵQ*�'7t��6"��ީv�����J�0` ��[R�2$7d��w��y�'!���R�����Y����2Q���^��oA�$���+�"�)���^a����G�ct0�����N�"���m�f��Ǜ�@Q�3�i��vf��O �J���UUJˤ%s���m�BK/*al����%����!�	� Et5;��Y0Jݙˏ�DM�C(��ЩKA@nq����z�+��C�����q��̩37Z��)	�&gZ�i՟����F�R���uE'�tʀ��`�"������ϓ4$��(�����vǽۅ��(��C����������AB��Ðq�V�A��^!�v.�!}D��U؟z�%2�4��w�-�;?�b����N����V���R�-�C�F�.��CO�xc��pm�0Ÿ�0%/��	D�\}�*���9�H�n]}�Ť�I��b$c>J�} �ۓj��y{UF>j�>��Ƨ#�e�}p1�>		�r��{��;Ɠ���U��y �.Ao*pZ���6":Z �xE�������]8��3	\��gι���H�/ą@�&�7)�g�v���R6f9! �����n9xƞ�Z��:�/}2�Ru��;z��7��Q������Vo���e���Q���m!��6 z�kw�]�)��<N�m8#�C��8��\r�m��{
{*�2��UnTܢV*�th�4�_(u�X�����l"������.���~"ֿ3�?=\��htg���6�0��_gd��["�k�0G2l}A�'Yw$��QyF���3tҌD� ���&M�i�#���u�p���� ��֥I�V�i#I�1��D���P����Kt6�h�sC����]��p��#cY����SBlѯ0�p���9��Gߎ#d<G�Bǚv��*�
׮��!o���<!�XZ�%w�b��Ҁ�2p�,C�hy�!Olt�S ���;��p	wSg�d���_�Y����+�{0��ѱ��Z������bc���2@�\�����K?��DWcBX�F��h\T�H��!����E�M�ȼ4�vv~ޢ����	�����h��Y���Ϫ	}����RE����a�t5l�n�Z���S_�C�`ʏ-�z�~@�v�҂4Lʬ�^���%��04�l����;��� �ݱ�΢�A��y�ze$-M6ޱ$i�Y*��]�%�yO���=	4�`��� ����W��dÌ���g3��=��K%f1���F���#�$�#6 ���tP~Pa��n���yڭ~�Z;�EbDGk�l�d���aB�\)�Dya|>l�+Ô#�R�� ������\Mj�=���}9ū���i�{�b���?����֮����Vs���4�Je�T�^�� ���9}�B� �?�#�I�/�Q>"����*��o'�{3I`�V�#�C3�0!��W�/�3B����$����VY���ֶ�eB]X���3|"_n	��O����I}�G�+�?/,�#�_ ��8󀘚�o��3ry;�,�-Gɵ@���Q�a��:l5"��8��O�RS.��	�$�q�	g�L�}-�xL1cb��,|I����Ҵ� ��w�w�0�����m��pg�O�R�	#��ktf�[���+-���C����������_d�p�b(����>_����"�c�l��ڴ݈<��
Lw�6U�������4ΉB���;�,�f�(_rA��Q}^wZ�K�O�A�<h9��5$�U���4(�aQ�3o[�Op�k��Y��`>��Ʈ##��n �a�n�� ����I�Pc	 �!�^Bڱ�uEg/:�m��S̗2�0��ou��g���]�w�Ñ��S�z���N�Ι�Y��*��KW&��tXX�W�<M�������U�͟_q��N�'�I��Uh��kr�Rz��z_SU2⵰p����p��>�7��${޶y˕֣��&���?�G��Üv��ǻ��-x��KטEֶ�N��jU�6��d6�"�v��e_�-ǗF�^nC���7!J��Jn�by!^�!������0��[��נ�]�s�`�;2����
��:��
���U��j�&�e��2�����dO�i,v6go^9��pkL%"�W}�Z���Aɍ��^����B���i�&i��&��M(B����>;m"
X9�Y�×z��µO�׊���^�[�,��k�p��!Lq��T��!t"�"cd>Q�?~�N�L��hF����M�ο�� ���.�0�ͫ��-M��*O�t��-!�}��4�v��03SD�*,�j� ��?˦�+�U��zW��EwB�w[��3�<ɏZ��?i*Tz�<`�0�96�;�Pp�S�)={��:p��\lP���x?8,��l���FB8qw��S���'��~P(��ծ,lI�5�<��7Q�^�"�b���LF��]��af��+���#u�� i�S���غK����[�!���Mzk��6�Zx!�� h���0�2�Z����Aհ���>���'׳��QF��2��>���*�2��?�rݲ�`�,��?���$���ju2����H0i�K�?e���M�O�TF�$�#)�n���i����h^�Y����I0D�aҕ�Ք�N �C\m��ˏՖ�N�F�\M�`R�n`�����x�+���K�[��hh�Y�ȁ��X�kW�F��j�[���~\l��qȖ@���� E��u�Ud�y-����(�\���p^��K���t���1b>B#PB�VZ
�Z�@%=�����v�����WLm�P��`Zrd {~��B��2 �G�r��߂�+�Q��/����3b�BQZ�n"J����X�h���|�)!6і}Ǿ�F������]�U�^.+�"�������n7Z���k�f(�?<��-�>}�@��"���RDx��:����P���(����x���V�l� &!��!�] b�*��\q2�����~��@9\�'͝xX �"r��T��"|2 k�x[��ips��Y�f�M� 8p�?�%XF��Y�2��uB�Z6��A�Ym�d�w�YP��4�/{����
��T���/����*$����F�>�C�

f��?Ŏ��V5r�g���̳�T�:+)h�v��GBR={�t��k���M������!܍��mT/h��W�ύ��`C ��,� l���d��7Ḑ&��:W ��g�;�מ�TQ'�Ȃ����G	���p<R\��EǙ	
��uq<elY�4`�������Am������60��L�{*���cޯ�?��֍�Ϋ�jS$�5z�O��/Qá,`�S��@�Q�{[Nb�JQb�m�_��X���x��4؅�[R����(�w�%��_8߅���_�����Pu��9P���_RR�Q���Z ��p�ޚX��yr:Qپ��ƶ��'gZ�����6@�nA��~��q�8 κ5m�3�w����)�w��l��gk�d�����١�^?U^���v������ީ��g��(��s������$���:|��[ٌ���3d8N1�]�4�3���~v�G��M�G�g���b��xHN$�<SU#��Q�2�cB�0��I�����������n.��:O[o��#��to.�S��Ү�G˞�=�a��ǆ�QV�!φK �ut^z�,�)���!&^���;��iI6y����u�Z-&���\z�Lq��kM��'
EIv&[5��x"#����Q[����*��%��:�A�d`3�6���.�!��>�[�C�I���S�����i����x\m�K��Q�B8w�7�7��#�2�f�J�(/2z��:ghJ�ԠSѧ�(>�3#��f׫��qS��J%��C��U�z=�֯݋Am�ǩ�ׇl�Q���W�q)Փ���LMI�s�0��2�\��J��F��+�"g�]�����@��o�	ܻ+��H��u�T:�M�b+�ǜ�BzR�R�T*�yK���b�ag�,F#$v�S�ù�Kɕ�<�lL�i^��0�o�]L��w��X��Q����3sY:����Ja��Fz�Q��N`*���[K�#���׺�n���3V`�TRkx�8�yf��ꌯ���ҧ��w��\�0���M�R�t�6���A��sx���È�I�n��G�?��ϸֵm%1N�������a��	�H��'V����#��iu�x���O�i�*�R[�0��J�#K�ʑU�4X8��ԛP�C%��� M!B�����<'��׫{ �v�μ)�ھ�%;d�=^+o�+^�����k���u�pX����k�{����蒮�	���W`�B+Gp.c�^�?ܱv*UGW�1ǧl^3��O�x���\�Dd�;��FǍ���h<��
�ĺm�v`(���T���mV>��1��g�ob����"ޤ@������l�iG����=�F��y����r��3���
�"����#��ؓ4�#��1���QU�#����^�O��M��q�Eb� ��c����[).N����.����kY���XKOӸ�P��e��6g�Ĭ����J�����9m�F�۷p%�����Ɇ���ċa�?�!+��B�1�R�|�Ӆ������$Q2���V�_d(�W�Y����OO1t��j�b��X���2vb�c�,�v(Cذ@��C���z�a��)�OM)�~o ��ֈ��az�+�t��1��d����|�Ib�r�A����W��<��e%B$�������zm�����x+��orl����IQ��B��N�	()Ǎz����ho��L�9B�i;�ި� ���9�	�8��v��E>x��3�?1r��b�_���΃�p5�fOz}Ne�ZX�� ��e�U��r�8x���E�:�-5�Nn�[ё�_
C��$$V�]���Rz~e�Ƃ��q��u���)��/���۽�7;\-*���g[e���wRM%@�a�0᧷�U��pKJ�:[��?6Q��Z�� ��p7;�,g]b�x�I9s�#��}��|����R�Nf�7Ѱ!(��� o9�8c@�!���T9ÉP�h�9I�i3x��Ym
��%�QG��ts�S���B����10Q��1l�%~1�Pod�`ٲ�x~�{��x����|*�+������/���ݥ�e�O�� �f�`�r&j�:�N�R�k+ٸ��Wc�&E��ؠ�wr�A.^4dw�Ip2̑K�r��<�,��>���c�w��-�i�F_�Qu�	2s�g�����۞r�#��ŧf���^K��1��K�Zc�DPz/9+�FӔy��t�_�E�F�`tf�J��8��!����Z����`+-�Jdz��)LG�Ơ]�"?هnp���zcU��d"�7*��]�WJ��P�q�,Q$��M��{"Z�4�2�,~��ö>M&K�e�Bٜ¯�ΧL]K�e�����8���DJ�c���<�<%0���Ι����Ғ�Ȝ9�+e]6�2��
�t/4��*�,Ug#���M�>��d�;��c䙖잽T�u�*��v�ݷ�5��p6�����W�T�{{�Q�]u���\3�����3}���C�yGA����x��Iؗ{p>�-�����B ݖ�d=��F�Y�jT��ge��$������M�&&]��[�N[C1��ײ²�,B���l�.��t�ə���o�p���<Q	��l#��[�10z	V(�aQlX��6��֕��`�g�D�_O[iڣ�̭�p	��x���mK�CE燺g�ky��[O��$qc��ͣ,���0�R���t�����,��e��c�m��)��s�	�*!�(��{!�d��=A��
!8�:��z=߹�����b�� ��d��[E���s�Ӑ|E'lU]]VD/T,P6�1,o��
��S��#_{�YZXոp��q_AJ��Yg�@� �(i�`���[_4�i$ϋT6�d[ =��!�Ϟ��I0Ϗ�HN]�@gu��b�uM�h}�[��x���95DRT�?'v���¿��a���Xʧ"x��R�)���-.0�"k`����n�����I�{�-��:X�-��r���׊7���­�	[�����S.�.ҟ��m�~���KX.Sk�i�T�ȵ���s�&%ʽW;$\��yIp2�xm&M>�F�w�GT����`�L�������َ%����7}Wy����p���9 �j���E�5�����V*j��2�&`^�N�b{���4�����%��'{\��e9neG*�c��_�/*�����S�¹��S���
k�<�7����z��Xs�ѯS Xϼ�:ơ:�̡�cLt�����*}��z9�OQ�;�n)(;<~�\�Z����=�ZSl����`�}�����E����8Eb�z�o�Z��9i��):@g'���[�qfQ�$ш��ђQ� )&0��ǧ�q^�����$C�g|�icl&�U�G��?�{U�����'
��f��P�=K�u&�U) � a�� ����a��yԒOJ*�����kFqlT��Z��;v&�E2ʃ���V��Z0�B�\9�������XI�D�Ȗ�Z��ƛ��g�"yq��z��W�:�y(.�jR�V����M��͐���W���2.b�����*J:���[-؉q��w
o��_������u��)e-��M��������v��n�g�F�s�?�ֹ��j�3=��H@"���6�'�(wn���H5fsW���4��z�n��Ʋmp�S��V���l�1�ؒ�z-ֿ4(p� 򂤸��M0�.X�@��
��?ٟ�`��R�JѢHu�������NC�/�Wfί�c�+\�+d���Q��"{_|��;Q��-�`�C+�D� l��:���-v_�cg:}7f��+:� �����6$T��۵��3�fK��4��s'I8���q(K��{�hV�]=Kl��J�	C1�Qk��ԧ�c�<���b�ֺzd2����J�Ⱥ#Z�����z�_X��.^��Y��� ��zF��Wa7�M��7��U�YS�yX~�uZ�\u$B����E�oF�m'�cG+O��,�2c9PS)�)��4�;���I��?���E�8��3^1bY� 1d����h\�?,���H�=q����-��k���ޭ=���n���^�,~hm���+3sMxz4��t��P4����%K�y L���`�>����X�����{���}��EK pB�~��x�3ʅ�#����Z��oM�Q�5�������Z#�5���(�Lg(��V����OsX�\�����u:�|�w]��՞��.u�2Tq�~��4MD��4;���Rh3^���,��C�.%F�#��	�6����:�%x(�+=��b 	��R^J��O|�9?ɾ�����cSB��tDNѱ���/��Y�����O%��	����r�� �h.��6�p���W:�~�}�nܡaU�����[^�g?7y�#�Ϗ͢cr��k���� U 􄈫0���B5$�k�}so��(a��>i��Z�O"��OR[���"q��&��X�Q���0s(B�b����|,?� 0K�=3(O#٪F��C�D�P���*��.j��W�d����t8�;sHT��5Q��"��FH�A�^I�ґ�M�Da@���'�xTuy_2�i�Q��-��P�o^���|4����՝�
�E[{���g(� �����J����Z� ����c��x��I�;(�d�0\1���",�J?�6á�� �{�&���St�[a�an�B�V\���*^ׄ���֒�֬]7��Ɵ �K��[&#F�&.��4��`��
2(���S��ij`�zAyG�3_�I�E�Ϫ�k��ȰR)�����R��Ӳv�Ag=[0���e
�8�#�x q	�Pe�bгϛ>�꽞tE$-ǃ"�DS�N|a��O��W0$z{�\"lÂr%� W�v?a3O\���� ����Ə�t=Ʊk@%��^F�Xuw��G��>޾�"��ٕ�j5�9J�F'kJ��� ��t�!u�LqG2�l�
�ȥ��@�yT��z�\�=כ~�+�@6<��r����V�?B�6˾��\�0�4��æ_�=�l���M#d�K<�������r����P�=�7�@��������/2Z^�^���c���.ō0���x�����K�H�8�Rk�����C/:.���
�쮫�@�c��Xk��1kJtM�&���$����~��w����1��t�'zO�{G�4R���E6#���V,"�ɺSl��ڳО�l�'d�UE�Ώ�,dIM�Y��	�*�'	p��cm�\� �8�N�ߍz�@\���o_�N%9��M\��w����=���)�@���%t��_&���5*���*�jd�y\Tk����x�<:�9b8Սq�dR �x�kī���F����FdTj&/�`'��O�LJ�HU]K8�(��&�K��9,����zrmv���xi8�
��yx��d߀��vX㫸�hp��V^sk�(=�S��̄v��f�j�z�#�0n�g_�M%���k��/�f�?���
��3jC�D�ӆg-�4�BY�u3ًa�꫐G�M�?4��V�z;*u�	����W���<�"�L���4H��}<l�cuu-9]�^��]�V�E�A�IS�� ��ʞ
j��\�a��x�%��<�50]�$[E�؍�+�²���_�J�beW?B��wp�����?�
��Vձ"�}�V"�~��Ӈ /�t�`@�%�[���)��t} OL9Yx�[��MZ�@fC������H�[��0 m/n֧�{p�+	r#]'}��f��Ø��0�����~�dZ�V����B��
�>G��.�1���?Ջ�)"���ֵi������f%�9�0\��w�Pc~n3we�F�w���2}�f��7E�g�d���%YT�ed�YE�)*��R����G�B+>"�:^�#/ L�C�F���@@���r��&�l�G/����m�{��Z�;�`�'�#�%!��c	X�ʭ�T�!��D�d/�;r��U2�J���O:2��ݥ��9$F�l4���wM�$���g\O���f�A5�ef	E�pj�T��;�����U���4�w�fY�.��x���>�\��c�ȉj����H ��&�f{�Lg�eE�yu롧m��b��N*AJ��M��!қ�Kf)}�<�]S��I�z����n�➺K�P��c�z�� ݱNcä��|Dj"Ļknҳ4W����x���4uWȂ�cNrgK����L�r��HK�U����}`�3J���b�$�z9��b���)���Nk��5[v�����|@�"���1J1b��쬌���Q�`Z��9�~ր5�H�>8��b-CY����BӢ^2��V۰�NWN���,��ɭ�u$�>(�,�nl�F�{�K��1
���t��p�z��� �kǭ�.,D�&G%Ϋ��V	�F�}�6�H���y~�5
>�k2D�8ʳt����}gh���v�6Ya���x���T����6mtZ��LXLpD/�׭���7�I?�8Ѥ1o Xm���S��+�� '��3���6�5�rg�Oč���RH*q�u)	a7o��X�j'�t�GW"U9:�|թ��.\�LS&�`��zo�^3�E9
$�%�p�z1�p�rO���U����_�Z;��D���򏺤3%��w�Ny8I�����-`�.�6����ș"$c�Q���Q[Z��7/�[4�k����v5��*X�	)���<�"ܗ���n�ވ��u)�����眨���>?걊f�IU��L��z��"�;��h�-���Ծ��H6�C�f�E%�sc��?*�6R=��bsl)��u�ODZ�m[�V�r^-���E�T4������.$��Б�WpA���'�\���	�a���%%��7��>vE�n�"�y"�X�[}hj�룷>�k�ڏ�wJ���%����S�'Pz���/���x	��PK��M!�%j08:��	W�e�qX#�G����p��4�����Q�`�א*_q�\ 6 |�b�9���U�r���L7��_P����Egdh�#<��g��S�OM�%,��a�א�'����"P�Ӕ�UBɇ���-�;n�o�B0��L���\u���H'��d��	�&�>�0c��:��s?6$��gQ���H>�V���R��vs��b\ۯ�?�B�hֵaL[���떔�>�l8r<6y�Є��΢��Bq��o��~�"�n9�./����z��\|X�D�d!�㌢A��"�����S'l�`x"׼S�N�'��X�J{��_�t��U�r"k$���B=w�y]�FF��\�,���1�Q�����!�y��L�߮K�01k_$V���D\@V<�&؃[bP,q��J���0���Y�p8���UU������Oթ�WW�\d��}´�}pl@�ޕڅ�7�u�ˎHV��	gl_8���i����H�q-ߝ��� )S�x �pO^g�Cu���W@��R�`"���vx���1T���Nn��w8��E&|<\�>M�a�Օe/��e`$���.G��փ��W�;̷�(��@�Ժx���3�ʅa�*�yȽ��F��/v�	�Ŧ��.�O�$!�?�E2"]�I_B{j��3�-,.X@���=O蚺_>j����O=�ő�������ޏ�zL�f���v�5�'�t.ԃ�}5�
���e��t�ӊ&��7��������(\G���1�o#:ǋ%PCab�Ȅ�z�Nʩ)��"���q�/8:2�ݼ����:�%A�۳���I���퀎��rF;,H��3�S���bn�٤�f��$���'�e�c�0��WH�"K��i#%�����ke�#Ke�	����:�k<C�c��P�0h��k!j�rZT�$��WM�eQ�<�,*�^�R�S锌��|CwW�i[=4fĒ($�������K�o����pn_D��j��ۿ��VüR/]�d}- �>6�7�`~�B�H�rk4�=�2���3;��B��ާ��qW����Kq��]k���6-::����;��7�h;[#
���TfN�5S%03�ǌ)e2��A�D���]�`e�B�@�hQ���Ҧ���z4�@�O�l�Jx���
�n�
}@�\O���B���YZ��ڰ�W�.68l[Q~
���K(�.M.^��q X���@;O��0Ϡ[}!�f� ����@1Ծej�����+�wE�A37
�A�?➰$��[n9���c,�^���;���۱ߵG�?�����6>f�Y���If�;���W�Ġ�`3=����i#4���T��g^�3�?�(}�T(��<��x2�8��zu��ʁ�m��<6Ӳ���B�����?�)�@�HJG��4��0���}f���p�k�߃]xO�h��q+י��EtC�>�nB��F34qR)��!y$d�:i�N48k���8Y�r����u��pq��w�kx`�-�ݏ힙F���): �E�5�UWkM6%)#sP������e��yHm��&Y�܃	��n[��,��J���X\.�%��3e����C�����!}L[`֯�F��N2�uN<G�x$Ȩh��.As�6��x��$�[4�EGu�|��ZN��,o5�m��ix���	Qwz�b���	��pڽ[DYA�8{*8�7�TA�tYz��q���ο.�>G��A�+z0\�Đ�>-v�RWX����ȷ�R�{<��T��J,ZX�nLbs.�~�
��Y�=Wu�������`δ~t�J#3��՗�x��_�z������b�v7��wC:��\i�HƓ
�|����%��!.Ǐ�1�?CU&�B��3T'�	����Ռrܠڬ+���F�^��ʁ�w�.�l;��噤?�3���1!?/w4A:�˸z�ny�$����-s�׊GpyYC0�U�gzܛ��u����ɧ�ݵ�vJ3Tk�Z ��6π��n�c����׌��*yS,'#�/3v��	�C;��Y��C�;G�w̽I%_#r�.�`��`�/Ԧ���Z��P�Mc���d�kX�.6{,΂�J1���	u���R}�s��&��G�`q�Vȸ�w�}�'=O�R�!yY��T2+�d�	V�T����[�;Ҧ
9xz�['��8s��gJ|--�U`�k^�����X�ӆ>��h� �^���-0�����1�?��3��x/��(K���y�������d��/�L6�d�ic��(#J�n��֢�lPv<�� ə
��z/A(��d]A6�у��Ruo�B��-݋R9`h�T�Ǵ��o�#���N,�2�H4��D*�M�잏��SE���ф"�Ъ�٠�@O޺����K���'�#[JÝLh��1!�E����U;6\��P�Ol�~K!�D��a�퇞R�|e���f���T���ҫ����k9�I�ɰ���Y�r�e���X[Qw��Q���:6k ]��ҙ#�["X�t���S?�ݡ���
��p3Omʥ��9��c,��hDP|�����g�����!�,�e���_�����t�n�,�J5���%P�|,�3�t���3�a��4"�����\��y�"���P����z͍,xHMC9Z�T�"h��r�h��X��&��f���]%�+�k�kS�,?�0��b. �Q(�G �(���@gX�0�1
Y�oy湺A6�nsq�l��ש��!?Fo��<ﵧ��R���me�Ѽ�(^������g�fxŹB���	�^���ƙS���藒A���KB�ՏR� E�)G�_��R3�? ���$=��b-�X�- Л������L�an��Ƣ����^� ���Z�c��L����Z��)o��m�{"t_pr�#nq b��.b���k��.@��(o�@���ߍ"e�4�[˳@�����T�F�T��@h�d��"�K7���o��ŧ��̓i|2�>Ԏan�4�˵>���Ε-�JEu�1Q���|��X��l����*miTQ6���\����S*����Vg~�����P:-y��t�y.��wԧE��kb�?�Pg�� ���U���,� �ld��_��詘�.*�R��[>5xakf��>%�}��8�!��-Q�y�x���+���u��ns;#��9�D&��c��wڰ�l���YE�P,�l����[�u���B�c�eL����z�~�13�J�rߒ&e�2z��J���Rsm�K�jT������ƙu2wx	i@@�G�]����k@|�$e
j��j��� �(��āɛi�h�cz�cqZ�Y���-�̉IȨ[^�\l�K�$�g�#{c��5·�Ң��iCc�X��2u���W���?)���x1D��/ ����+]�0q\Fл�,Jx�������W��r��昷��r,L�f�F�.��
k��C%���
۟��?�Nm�O9�4珩1%������OUP�����CG��6��gYjs�������Z���ϊOA�t��$�nD�1�o���"Ԛ�Ĵ���G�l7���4/�}ٛ����v(���W��BW&�훯�����e �39�ߪ@�ؠ\c~���Σ���(ry����^�*=�rߌ�_� I"����Ŕ��!V��ƽ�Ȃ�p���G�
]�My�#,�ޤ���k�G^�B���H~�Fa�"^Q��H�����(YE�	���"����5:���)�>��\��Z��N���{�:�U+L����Z{����N
�Duù�x��L��M|Sd�:�(�5��jZ�>fa6N�X�G��-�����k�Q�M���,�0���G�� �֏�q�.~��o�_B̽���B��)�HSE� n��`��v�Q�C.�[#��^V��-a�F����9^ݘ�1�L�G���>���y�*����E��ΓOy<3mDj�E�0c>��1~H�@y𩺹�aipAC�Vл�3��ګ|����H��K>yv�O��n��3K����2w�3rS��V��f ��5��I�0/��� �H�ՙBFJ��m��$�d�շ�!O��BI�}����:���`
!Q�^�Fn�3vo��3Z��v2|p�7>��b�l����L&^t{�0���+��x�����44���:B�JԶT��)���ҋŢ�-�ķ��ؽDM�<05ܕ�F��!h��y��c�$�/+Y�e�a������,l��k��CyV,�@� rZ�I��K�0+u�|<Q>��1+37:<�:J�S��5��|!-���yW�)����L���Ǚo�<��L��%,�p�8���L!�6�(�\����rϢ�6w@Ev_��K��'!NB%P���\U'����B�`�9��O	�;=jQ��d�S^�VK&Fl�T5�Q��h�����\IK7ֿ� .=S�������]�YMҺ�WCSp`�]�"T��ͣ�����j�l*.*��Wߘ�+u����P��w%\b����}@\�߃՜�����?WT���"0񙹼��Ģ�i\&Q�����Ԕ;f|?�xU������$N�A��_�����% ��9�����������uy�A�[�b�CL`���5�(#w�9}'�Ū7�����D�Z_�,'P3!�$�H��,x�L��i��$�4\^����Qt�t��o�[g�ݯ�寇	�ޔГIb�ny�2��0"I� ��vD�'=��(jc9K�Ϣf)���P��e��{H�Ґ��G�۰�����&+F�_<s�*c;�0*���Y1�dk_{�a]�^�j���Q���z�ӨE�:����C���o��~��^eW�=y�~D�Y�-��\�O%߆j]?��`�5{!q��d M��J5���>O��.P�?�sU������X>�+e�@����5-���+oG	ɕ��i�wP:*�5�N��|������(��l���/��?��Jt��g@ &�Y�ͺ�Z�E�،i�?K�朴v":˗����mǗf(���$� fmp����ؠ�n ��z/��A^I��I�����\vQ���I�$��Շ[`8�Xh�����^�Z<%LX�r�%�'�����ASp����k�kk�7 �p�j�5OX)<g�\���-9��.9)����-B��X��/�bG��%�=}�ΑVmco��涎(\m�Ǵ�h`��d�}�[��d�E��<�g��b��0o�/��CJa/�e��pU�Ed��I!�M����U�-e��S�3_]���O2�|��Y�59��s�<J%N캌���1�Wby�����PH;x����qXd�B�p� !G�H�F�y[ƾw�u"2���=���e����P��X��8Y��ɺXꈛ���(/\(�;8]�:R����\��)���������f�.�P�?Wc[tW8׫)d���܉q8n���P�5��9�2h���x�9-�"B}�� J?sl�����(�V��Ȝ���	�f�X_$���x��b�G���`)�a>��{��Z�vT�z�2HE����(��- {N��.�õ�p,\�������IJ���5�C6���X#\O %_\�UpC��6k��d	�7��RL�5ӆ��;p���~i�1��E5�a�b�����}Oc�)`&���R�8;�D3�!���-W�����L�
�H�ѡ��6��TQ(S�>���@fz&���j�-�~z�i�ħvmL��&�EZ
>h�gWܞ�#�xm}�{'d��ع}����AV��;/.ǖ���Z.�-\�K����K��))�l=+��g�	�no������m���R�'>�B�"f��֗����OZ.Oy�5����f���͆��g�)�ʸ��H���b�\f��~ڶ��A{��4ɦ�|��yG�t�-4�ϡ���U޹����n4�J4��D�3��� ���iN7r�᪫�eQ�Z
ao���������@��n��n�� #q�Q�j�}I��>�XiX�0x۔��-_w0�Έ�����h��Z���	2�1M�`�p�:�j�a�nD��
8���C*���?�$�萢x
���(�
��{:Qӟ����v!W�*��������{j�Ų�k`�vX�V䩂�T|��&nT��*�C�.��zgɞ���T'@��@Ψ�~0�sn�g���Ӂ�6���F�
93�8ƴ��Pl� �$<@��gq�eOK�υ�&w�քu}'�x���H~Cʜ�z�l�����^��B�q"���C2���#�C:����eĞu���rH u�U����YU�Y�J����mQJ	��^��:��	��S��M���W�Q�Kf�P��4B��^֚Zfzno�)��.n�)q�H�To�/g(I�<�D��Ulk�6��2M�3��������se��������:�@�26�z$9m��!J���r��b���/��m~�nO�NX�s]~����k�������QK�7��a���?�w��/�Bp�>�y�)0ۨ}��F�DB<I�R�k����on_LL�Y�I)w�*չ��N����@��Ui�C�UĞ!�k=K�]q��a#�e�Y����oĮD2���R=���}�~�&H���SP܅VJ���U�93���'�*J�w"j
h4c�h���[�F���G��=fYt+w/��UT��`πC�Yn[g���L�-7>V�o��|LAg�nVLKmTsz�De��u'�]��)�6]�-���D���I0��%zk�	Qe������+���e+:^��KKp3Z�ĬQ�e���Ie�eƍ�*'~�¦%2�T�h/�u��ob���t���}��Kf[�hl���P TS.bi ��W �����]���`��,-Y�ꔃE���Ǒ�hY�f53)6���"92�����BOJ�G��</3����#�O{T&�c�,�'Zmx��Ϟ4�����h�~*U��.��D{��N�ml�v��s���C���\X�rE�ED#�zՔ\OXJ
B��3iF����S���j� �4z�j�V���\C�91��>Û-�"�%ϸ��yw:n�~����B�+]�U�2s|6�^�9G�͂����h������_Y� �Ncb�S�w0�Tw��6W� ��MsU+�C6��������n�4���Z?��J���Tm(l�GŐi6G����1�zvZa������zb^'���^��B'��Y���P��ri/�xЁWT�9�jw�
�ӌk&�6קij�<�zp6�M�#�K�lx�74~=?E����z۴3���	8�j�A4��&4�].D|�m�
��}B�l�)�7�?��M�L�+�_A ��Ҵ�$�)�������}�5C�vBf#ZKaOp�C�y��絗x� �Q�t���ˠ���nWR�g2��a �'�P��9<�5�R��>v��?��aՠd�&��.�7Pc�q���X��Elb-� ��_��v�������mj��q2^K�`^���nJa�x�	 �И�j0�k�r�q�unH�d���3�Ԟ×G\Ow(�$�]S������^�}^�t�wK��Pz?9ߦ,��hS�c �1��#fp��ݷ��b!�V�����Ta(��-$4@e��g��P�Jg�݈?M��F)H����lr�B� ��pT"����b�}����/���@�f׍ԑW�jqK���oҺR�s���T����<�U!v𖢧Ԃ��Wކ\汘�E,����[�IU8|��S1�Gc�=ׂolY�H�/�(�E�����r��pZ��2L\�V���EC��TJ2�rJ`C
FOɠIN��|�7OB��<�[�$b^��i��tY*��ϝ��$�ukF���Z��W�:Y����h��~�襞�	Q=�q�P�妜	l0U�S'Ǡ�➸lI����B��(�K��Ҭjr��LK{g?���ZA�4K��b����7����[���n�K���DA�Q@�ػc+V���G&��9�hh,��'��ƩO�V0�§wGU��l7ZU�Ȁ!�i0����H�jZM�La`���*,��@��3��v�Ni�n�N��6�A.'	'��۴:KKU�|K�t(<�D4H R�u��>�5I�-Ų����w54�����M�z����ɜ�PK��6���~��%7s�Q�s*Ϊ�x���8gw�[��1A���ޜ	J�2\��H~�߰@���od˙T�^MV����_sKJ�)ߩO��a��7)e/SAV���A-	+���e>��H�hkk�1�]x����8KJ��NRg]�15w0/�	���s�o}4r���B �E!��fJ�-�8(2��-!>�,���V"Ѭ%\w{3	�0쓙b�6�X�#�=��l?ko[�.Z���N��B�j�6�
�mO�Sۼۙ���Q�@���0�8��苝hYp��,�+��q�c�&-}�
��ԅ89d�t��Lw���7a��*��}�+;�㨖>�[(]:A���Ȃ�s���S��pg�����<4��w��53劓d�T��A�Ȋ}m������!�U�+��yl2=�kҟl�!o+V����o3Jᵮ+4�J�f;ڷ�&L�W��RCѲ�F��-��֎8�ך#c��R�ʞG"j�N���O v�M���O�d�L�g���?c�l4���*���j�-y�A�d@V)P�����c�'O���y/������|Ǿ� �Mj���|��u ��M���9�>!�I�XI緘w1lhwެ�BgF��I���%V�ǝ/|�jƪ��165�Pح��dS�9�ᷡ��w3u��ɬ����n+o����=���ڡl�ּ��Xf�6߭����"���{^a��"��m0%<�v��n�ܬ�	��(d�ijT���>8EE�ZSw�GA�7�����)��o��񑒅A"��j��xMf��֬�$������"V&^@`a.T��Ւ��?KԋMY���A�����;z �!$w"6I: ��2���<ʷ3ۨ� ���֘�|��As�!�;d�ʈR.���Y�Q�4�ǧ/�*�y��*V��.�l-aw*"���;A�����P4DScU�4��Zg⸗�s�{O���LP���[��̱�>��c���o �̱�����ۦ~�1��.m���r�q��{�gaʇ�I����g����u�rcS�����ڽ1#��挛Oh�h�Z!;G��#K4�!¸�#5�;����I0��5����z�q`�݊���4�`4!��mP�����_��덦� ��.tPT<�� p���tF^EEd�i]�Q�N������wE2�9�aO��R-8S��Z)\k�fv�g������k��y�&�6�͑	��o��'�V��0=M,�
����R;P��� hs�����Ϯ�<��#�XH��,;*�|�RG�o��s~R'I4�7���������S�L���G�����H7��%��d��g7���
ڜG�����G_�v~^+
�^��B���,A0�?NRz/��Ȱ��i�u��,�FUA������-��%�>]�r�G�b�mx�k`��M�1d�8֎�.WL1J��} q�'�K�h��b�|����z���UQ���s��&O���/�v%�5wme���]�gYW�;,V?�V�eO��1�Z�O���*ez�ВT���
g�,J	<|n�4�o�:1�I��Z�Y>�Z�j�/��#--*�N+K��D]$�Z�D�euN�AA��q�/�Tn��ڲ �D�R����ħm��|�V�vVC0�;�?��ܧ��w�[<Pp�8w̛".,��/�1K�G���P�eFN�����]�'�S�w�i��r�܇���ع�v�;�ט^gD�X�3MR��`N^�Kwa^�{����d��c0z���{�I~z�}0��щh�����ٯ}Π��|�v_�,:�_Ah�� ���F"��ڐ�����ǀ�ׂ}e#Ծިbl���"�ۑ�J�Z�!VCZ1��FC�n�!�I7�4�h�X���uټ!���>���.MѤn+����z����ғ&���+�I{}c���}(}�t�W߄�b|��}Q���_�M.��;�ļ���ǚ(^���`�#�z_Ke�}KAɄ�Z�j4����K���=�F�1��:
����p����|���8��s��ly���!��ݳZ6R,Z�c��5Y8�U���g�i|ar)l��%S�owi�gm��Ct�t�䄒��B+x��DW��3�g�,cJ8 ǽ��T�h�3Whj����i���C&J��Q�ұR�i�?X1�qS���Bv����QU�-��{[,�ʟ��oD+���R�u	���ņI�G��&f�2NdИ�ۏ��{���3v��]D����8ի���D>}�Ȓ;�WJu���CO��^�6��%&8^�Z���ë�h�f%n{�;(����5!)%����M���1�ّ|���g���l�8K��8�3��{
�#�� ��c� �A,����3i-����	��VS��=���!tR�Ŝ)���"�<��#��ѲmD'fn�\�aw��:=�=o�ƀ�ai�\���4$#	xb����A��ӕD�Y�x�ß�
��2�ŠSs��j{]���g�(*�m%��}Q��A&��o>ϧ_
�R��!"���(�Z�*QQxi	U��/M*�N��Y��Fn_��L&JiҮ۱I�3[���1����L��*�����RJb
u������t���2z��<~�,%Cb#1�ϩ�T��i�b.���Mq�_��~�[ߔG�ڄ8Q�-*3h2��_i��P�����;��s��&�H\k�f�E|Cei��6"P��VB^"0P@�;���1&79��s�ǋ[^����k�M���	,4��A�rEQ[Ǩo�/�ς� �TbG����s��|�7�`��D�N�L�� �s��K�Ec�$~@���u��}�)���#wd��5�L���M���&�?��!y�sDT�`�v3��}|�dVe�Z�PX=r2d�O�r��v���_7�{��#Z�`O���~�j!��1B�48f��ax��d�ȇ���sp���j��w���f�\(dm��p��l��W��= �:ƝG�h�vR��z���钭�=ƒ�ג7xZƌ��4�WDU�Nb�~�9>�U?����%	ӧ�G�X.�ƽb�I�iM������n�s?ǚ�Y��������C3f��v��=�۝Z�������E8Y�z��Zp|;���;����� ��r�ݐ�?���as�;�ضe���6
0�:In�Y��f9��F�L(������NI&�'��D;t,��L�PsL$�pL�	L_� X�.H��" �x '�~�-��h;дau��M����Ϗ�b�ȹζ�g,�2_��U����i�-��`.��گYY4kX��p;�2����k�w�����H$��4�<{�Km�&�,����m�.�q��ó>X}�h�y �������	�������#!9��$sCy�o�N��0���c��\�A�w4��a��1"}����uJ�s0���3N5�d�w�q6���or��PE�"��#j[ŰL�!�@Xٚ(�q� cz��p�I���.>��eՈ���V��W�c�9p��� Y�v����\�㫕Nb����.�xE����,(CK�}g�*�
P߽�4�=��<�̳��WT̵U�������óu��P�P岁+	�1�R��J��U��;*�st-�e����Љ��СDUU�3����0�k7��������;)��(�1V�?�4�~8�ƽ ���^k�5K���^�Y	8��a���C��=wx>�rwva4���Ө{��:��Ӹuss�V��gu2K��7�4�0{���f:w2�^�{�Kt�U���=��F!��^��lq�M۹�����hLb�4��Ի�ɿ���6r۽�#�z>�a�,����0�7�댐�W���X��bz�e�F��Ul�o~Ĵ�.�A9�MZw��vv�[&5��c�:6ɔ"^�Ӣ-!�d����S�6!i��f$*��?_H⼈���p��rK�~�g3|���U`p/v��]�Z�ܳPP�)�pUƢ�������&D"������)y����{w
�1:8.<6����{�,�	�9�Ֆ���ѹ�X!���"i���{��7�,^��u���p�����lj}c��
`�/������]_�������9�ķ��q8�6Lذ�	1�T_9��7.�("W�庄����sD�ڤ��)�0�+�K���۳�/�Z����( s3��]��xA���/��#@O�	�U�:l`L��Dh��"�>B���3��{3H�ɯ��[��۴���V��5@��1�V�T�L�^X���sTlť%��?�n��عqQ,�J��g��Y��G)�8+^�K�[�>{P�.:P���'ߖb(�'�2-��n�P^��K4����&�������c����YV��ݽ9� �&�П����{��@MA��X`g�
e���c���P�T�z�~p�H�F5U��*:��8�WЛ{J@F��9-���O��7�+z��$�6�Qc�b� ��ծm�h/2�3���+�p���=ƻU/A�v��:���~���	S�����}��'6&�T<gPv'	8��P��·��S*"nh^iJ�����&!i �:��l����+Ð�������	��@d��팇m�1o�YcQ6^��Ǡ���{���~x��՘i��vI��hn %��t���(,�ǳ�^�G=!��~?Q��v�^B����c���;���_~P���2/�1�)��Ƚ����&Vm�-��)@u��9��S��p�8��б��L�����P��e�C���V�8-ᘶa���tEevd���E��.�@�Tg��N��@
@6��l>Y�y�~�^H�Y��]�vwtЊצ۟��r}j7�-Ȁޟ���d~���ĿՁ�㺌0�[=�G閟S�:Yw����j<c:��9<[�I�Ѫ��c���R)��S;��_�d<�b6�:P
�j��*.l�zz&,���?�=�~G�-��G��	B	���E��R6G�Q�T�_���|S�X'�u�.p..]����������
b=oG8��;��JfLP�k��,9��(�P3U������Z�W*��4��"���8� ߸����?���G��`�I�̿�?=Z���`�kU���56�3.��B�n$�Ѯ�Ӵ��|.�*���L��$�lV��ܮ���'.L�)|��|�����"7z#�!x�,���q��h��KBU�鵱��-�H��r�\>�2q��1�z���g�<�mD�[�]��.3n�1ʷ8��M�?lwQ�X�uwX	��?U[�\X�G;�gb��u��t	_��!9�)�����+Q��
�����d"н̖Ko.Q)�z2&�͊�_�D#��~�?�>��+E���7
����65vL���&��]��-��Ǆ������'� 4+��@�����qx�
3J�j���އ58:|��z���s���d�� }ԯ���òM:	�7�U�:{=h� d�a ?=�"fD��F�?�ژ��餚$�mujl�.���.%V����rN\1�.�M�`�0��\cu��1��p:X�n��[af�ձH/�P�1��Tʱ����!�n�+�54�S\��MX���¢6Xr O}�}�����T�0���BO�_n���;kp�I�%[��@�Z#_-��ʀ̡��Ld^�����H���⫪�u��� ���{�?hab���H�����rO���/��B?!P����P��c�9�����gI�����R?���K�S��JN�2���p��՗q�N,�^�Ͻ	�����I�)m6�^i�k�Ohdǋ��-��'�c��νB =4'��LM�%D��y\��V�$��l�ΘFB���D4����Da�H=��P{��s�.�Ę�����g6e�ҧ��MC!�7�@m��&7,f�}8w�'!6�����ӏ�l�&~vƬ��O��>����&֎�1�DB�p�£�����qɟ��.N���5"��-=K�J�KB� �$==���D����6�X�}\�M��=���l�<V���**�(���K����p����㶶��
��U=B�����<S�Mؓ�dt��[3�q\���� U�!�[&i#FUc��ݔqX|��녍��PP��N�a@�v���V�^|Mu9�ޛs`Z�E��v�Zͱ��};��In�_�a���8k�؏'-��ٷkE:��\�Q��G�϶�+���*e%��������$J��çiތ[����A�������'R*���]��/�3NjK@/Nv�X���p�*k9�(���!�D����D�h�Q�o���%D�?;�hf4$	!��MP����#b�m��_H�y������S����eG ZMWjJ�9���'�ra����w˙.=n�{��7>ƅ pQ�K�
���h�څm,�Et���ҏ[�����K�&�����j>�ZՅ�t�>����M�svɞ�� }��������s/���;���;���c����@of�.��0��xe��ȱ
,J��[��|T�]2��n���(���rG5�2���D��Gǲ�<�	�?g\bJ*n�q�!�6�����ң�����$�8��O&�'�H/ir�v̜�|y �ufާl�l�٭�zƷ"`�O�7*V��xų�*F�I�뤼��Q�``�^"�Q��&[���e�����#p���ۈ�C>�b��oB��*?���ӂ�V8Av$ 5Dj�B����$<����I9��S����=�{���Ҳ�b�$����᝞��z��=��#"+lK�j�z�ȷIG��������> M��t����a�D~�F#��aa.��Y殥B�Y������ k�"ZÑ̰����Z�S��q��B��ct���Q�>1S^{�/��{a3�u<���1�ޞe*#([Ed�%�rCK1U�f(���+ �\'��W�Z�L����ӛg�2!�aU�p��T(A�����c��<c����eG�d���y:X�P�@]�_�����gM9F�yg�LړZ0���Z���r�����p�����F��洎I���+ O�:�H�=�~�J���c,xS.�tB'�6�]F��m��������S��Y�9m��L~�r�L�̷pf�MP�^{�|m�u��<��6�᬴�L]�gC����p�NS_ۇ�$z ���5�o��6!L�d��|�R0�֟a�m�h�T�G��Xdh� /.(���	��&��RA̡@�;��eˑ$ٗ}�7��Z-�3��k����Y��9k�t�ȗemq_�"{/�n�sfB����i�(Ǒh���o�q��I�kS ��������Iߎ/��N^�H��Z�貶G	@;�m6קs���E��*줢�,[[+�����%8V1�&1��gD4�C&�!V{�<ה�	�吧8����K��/�m�m�LO.��|[�����Jp�y_jz�[���Z�|�R����Z��FUAL�4��
XS�Lp��'N�Bhͦ�(�Ƌ�I4-=k��V)���G)&�a/J��1z��E��U$t>���;������j�aEܸ]��R9M'�|Yz�S��7j4v�C�	�$�~�5����دx�g�*mQ�����P�p�u!;���݉iH�+~��%�\Cg��qZq_ˢ"�d�:Z&�v)"�u���:s���h�f�o>��N�v��s
���oWo�О?M3�~�@���+{�V�4Y1�,M�l�ˬ)-I�X��#m֩ab��Ő�����Ɨ������}�a�z����fQe��+'`Q��;d0�ߩH�n�<>��h��`�\���6�T��n�z�(P�n�B�`pt�7����@|�ȥ� J��e͒z��ؠ��=��pܟ��JdddnH�,�:�u�Gn��:�Zf���	e�����uJ7s�O���x'�	,Ë1o��^;���$�#���$V�^g1���y�&�������}$Nv��q����;��E���o�G�m,K��u��z(p�� r	57|I¡��Ѓ��3���a�m�HW9�N��)���Y
^,�u� =�d�74*�����l�W�`��E�~;�������p�@��*Yr̕w��@��렸��݄�^��r`vZ��r�����_�]��E�`_��z�Rz�B�Nݾ�/�t��(��iS6�g�`ꭞ��5�RG᱄�	�3���J�� � N�[�c
�2�u�R�[ �o���M5��9j���$"K��l�~�6%���RL��ʗoJ��v���vaZ	=��$Z��gFQ��*�d�7B��Il:�K���>���@,-(��&g�&{���9�*#�8G]�'z��*n�O���n����,�E\.*Y>���DC'���W�3l��&	�=KR��x�����4�&��.H�Sl}+A��eN��~�'7	/W.���?�Py���A�WwPq%2[5:���g�;�� u�C ��h�Ad����j��``.{�ό�WF>}=ͬ%:Z� )��e.�3���R����Q\׶;�:�����޵D���#(7�a�6��X�3��K��qa�7�r�w��Ҟ����(�z�i�n,�F� ��2�I�x@Z���_���fKߑuI�>jK�L����ͨ>�6�x������g��"5��B��Q��9��Y�u�W|�)5?����]PNS�8��� p��z�]a)�w�RTW��ǿ�q��e=RU9!�KX2�[��_]1�ʐ��I�y-���U]m�=��V��?�"��m{ܿ·��J�Bw�,�2ײM��I{cl�-��q�23�M��;�R7sb�w���c�/�m0�0��^�!Џؐ��K���a���l���Ȝ�J^P��� ���1�u	�?��b4�A��HP[e8�ep:�*+�Y-KO�?%jC�B����l���:7�9�>�ջ��g{�O{�ъ���|�-;��+��y�'DgT����Az9�ԅ�����*��|�,hy�E� ��XKibºO�y*)�N"?���l�g��n����v(
{k���n��瀊W)���M����}�G�J�)�l���{��SM9�hJ��D�xF�fkP_�r��i:d�F�;0�z.{'6�C�r��ץ6l�J��pA8])���m��Bkk������r�F�8
/�`O&Ʊ��[B���K�b*�$$�����wv�cs�ڕ{=�V�Dr��4�v�U=�TUY�x$d���͆��u�^�k~Dz��*��^�&p1R�җ�E���D�%�P��`X����2i���X��t�Ny�jcf8�kGp�u\���cX�)���n�xM�:�b�)d�eӽ�^i't�ѫ�<L4MF�W?��!��jυ�":S�U����u?,��q���)�V� }Z��&��VGɭz/E@��YN�rX���3���q�7u�=m�٬DUv���]Y��Z
��o��lD5��fw*N�kZ��i����b�8
�\�"ϲ�`��=ܐ�v��,[�fc|�;1��ݩDL��Uě��Do5@��i��`�(��B�-/ﳆ��f�K�]���2�ʸޭ�����$�`
�nr�(f�i�{��mS����, /��C;/Ы" s�w�m��I+T���5UK̭ V�
n0\T�^�Z��U�P���3��FJzD"���0��we|���
k�P����e����g& jC�+��s,Tsc/U��v�5U���P{g��Cr(-�7�2]�0�g�L'U(�}��Ҿhm
t �_�B�V2ʋ�<{����G��>:7[�T�qB	��� �]���^۬Wy�9 x(��DE]h��>��6��l*t<�J9��ߪ;\Tm���`����o�S�:�,Eފl��tm�۷c�n��i�SP$D7��������C���������5f��r��.�|���aNtWU�뼃��:á��P����c���vܧF�=<$�tYMhqd{k�Ӟ�lDA|��l�Q�_��2I�eXW~�{f$��Du�!#��5�jyh�sW+l��F��I2�.is���)t<T>$@a`��K��2! ���`��ʧ� �1��oX�MB"}9)�w����*��d0a�7����U�x4�h>��&&O�4�e��\��`Ց? Q�y����Z�f����������B|��>x�-��5������E�j���bB�pq���B� `�C��� ���$9���;�|PG`��S?je��d�82�*8�<_���
��O�9�4�V��wnz�W�Fb�"�@�&߆�z�'!�ePq�s
���R�ޞ�<`�����b33�.��������2�}
G�~j������n���:�qS���ګ��(�$�<B�_�?�X8 W�^<�wWz{��/t�Wc��B����m�f8]��1G�]Jۮ��U|�����K��jõǑY���w](T���w`�OKo�̐TZe�CaEb;%M���;�Ck�Qk��<�����9g��
�\qt(\0^���,�+j�uC�#T?�șL8��0��Ґ5�AE��]<]H�,:A�V� ��� �i�t��vP  %�I?�����f�Js�-�w|�<�*�%y���g��3҅��\�4Z�DC�-z�v3\f3j-�iU>62��?�E��w����d�u�M���{��E�� �U&�@����}ە�#Cl����x�:I`se�%�\I��y'��Ƒ�c��xÐO-z�y&8�k0$.3���$Z��W�p)O�d�6}�2U�->u)��qζ��Cr�\AW�İ���˩_���0��pO��z'��M��!�,��焑^a��p��fK�3��-�AyY�%M�	"k����6�YʌY=\,�z@RR_֦Xn���!��\ûSD����w"�W���=�ko��5�?����Ϭ�|��ļ9��}�T&����AIpq䨐	�J@ ���Mm@ ח�^������\����4[ZO�$��<ťH�ㅚ`
���=#҇1����L]�Rw���~�>���+�d�A�����{�che}�Q�	~�g�~� �٫�}AI�WWVW�@U9�����Ჾ���6��5�.��B�1�C�=�1�c��L����4�{�0�!$�=� Y�,EM���NՠxG��Ps�:�?��Vv{T�k��a\��Du�#>=��������G�}�������8A"X	۝�#�N�,R���^\�洽����D*��Ҩ����4��wV���c����m�u�eE�t]A����=���XUe�y�	�Z�Y�r	���P��=���2�����mm/����*�-.�.�]��Sy�i��{�*:�m]M�ð;\�J�ٷ�G-������KL��^��MDB��źV=��v^���,��hI̞���*H5�gt���7i�Tω|+�E/����\J����5�cX�7���J�عIKH���/v�B��Ծ�P���*��s������?���MԾ���u��$|����3TpBS��謎���Pƕ��2�2�~Ɵ
��
"U�76ZW���Ooj��?o�(#宱��m�+���BL�&v�EJr �����9�`惔"&-��[���2����xF�:�!�'oP���eݕ��
?(t��^�䎑�>���t�LӳlT���D� n��4',wJ͒p���DJ]�r��8F?=Nf�wBv��>@�p��?i�*x���|�|�?6f^w�Gz���M��
� �b�6;F�8ь_r~m�hq�JǠc����)�7��4î��I�k�,���^�j���ՁF��c��ձ�	2��;��qE\�_�eT_Q�Z���n�!����y�.q;��F�@���9o1c��Q��R���W����"$؃�Z,˪b�f�Oȶ��-�V��K�k�s�oA���Ԉ�s/�D�8�qT-^ZE�@Z��8ϴ�o>׃W�d�KX�3oQyQn�]
����q��Ї0w��NL�k��=�J�<��9H�%��9�
�܅�dTp��zf�,	22(hW�+��!�W�V�{of
�55�z��@��'�&�q��:��'�&�;��u���e"3CiOW z�<\P4\}�v�Μw\��/<��p��1Wo����bK� �M%lȨ�JSy_䜜��V����R���z:�^aZ|��3��Zxyfj����E 	��"����`�'�v ���N6ghW�s�\3Okoo��)�Q!L����2Ū��O��U���8V0���w��
�I�]���Y]�8(����]�ML`5�#77|�2=C�O��!��{g�}��`���]��l<~(*Z���+V�|�Ӵ�*H�&�%�v^�m�E,��ay�K{"��u�����o�Y6��Fc�����
rq�g��s��uF.凯�T�����hjm���T J�XJ�̚A�)u�����Ӆ������4X���E9i�����vq�M�+R�5cl�*!��0>��aL����I���q8H���	�a�Ik�\�?_��U�(6�Ǿ���`� ?�Ҙ��(���3�#�+ZQƎ�ttl�^�}�:Ɛ�̸�Ɉ�UI:���E��Q0�H.�*��AK��?ɖ(o���lO��������XH�7!��im���t��.7V@b^p�;L�-�Sz#Wl�ة���y��>�1��v%3�J�3�ɵ$�`�����9u$��2N*�O����rnf\2���q��������mxH�w�����UU!��Ͱg���5�m��偎�1�|�?���0C ��h�X"��Y!��|8NGT��O�󿌁�DP��B��Dk&�X���#e\�!�� e+�9��Vb5�1o��Q���-��`�y�dΠ����)8��-��Ѕ���.�[�*��g��9�6�_�x��b��(�r��GԿ
/�z����X�}��OЭ�%��s�<7EZ4�C�U�Um�C�	�b6��`��,�t(��][�a�K:�I=��|�(:vTW3��m���@�JC�u��deU�#]��#Rf��mz�0�a#�I�ʃg~�,����F���\����&|�쳢Os���:�]~f̀wx�D��yG��ܿ@,�?1,�Ŧa4?�̟�[cwѡ$au������[�޸�rO��W�sU}F��UHp�y����%��z�S-��z���[�`�}��b��B0���v�r�E�m���FYf���%Ad)w�+�^�Q��,�:��N�.�>�G}2Xdq_�!(�N�Q̜�����U������ܬ�t����:#�ñX׮Jdwg/I�����U��W�M`�w]b|��@EP[F��P��)�>E�	&�f��4K�����e�@����X�S@(v|�"��]���+�$�Wm����a���ވc�j��OsY(1.d�ľ
idic�L'�HH��cp��1W <���$������ݓ�̄yA,�I�ѧh�����y����H;eҐ�=S�����g�k1>S�ٮ�¨31�P�|�[��f+X���Os�q��!��蕢����������bg��3|Y�wO���(�$��#���S��LK�Q]6�7�Gv���"�>E'���Ӯd��;w��'Ɂ(^b���k�����+��t��[d�`�,�Q7�g)=�����k�Q����	β�ba�uc�b!�bzJ�5ǞX�R���jk%S��c^H;�
`��2�g` �ԂCMh��-����y�Q�zP83�\e(�1h�K�a|M�jY�)a�T6�9�	+h����CՈb
�[���k�O_Bjf�)HRC$�������hI��
������k���1���r�=P<F�4+&�vO����"2Ч�C���_�t�ઔ�Pa��}L��,e ��)�>-C�ge��%s��S� ��r��E�zp���e�pZ��v�X�ev3G�{�%Ca��?�?c5�&Q��J)'��O�5�
MM���-���KO)��rSh�*��?�1�!��3�:�N!���Hq���զ9�%�uZ?$\����A�d���|���g� ��dD�����5X�ژ�;��T�-�Lib��r�i"jqe�=��x����M��׽���Z�0+Gy�<3O����ZN����U2���P~��62�A��'�~���qɆ༓x�H
�r�{� ��oa�[�Է:�$�	hM����ý
�2��Rd���={shu����̖���7�#�r��@=�3J�@���r7�ݬ��ٗU�W�dDɻ��`;OTIze��=�ml�]�L]\�\�SX'͘h���
Y_g��_F�'&������Ң~tvRt?�NQ���������Hi1��0 ֦7/`s��W�D�9���%�໏kA��tM���^ץ�>Y�]��d�oT�N䅓L-�WIw���!��)���I*��������M�'=�v�Zb��n�@?}���o�QϪ 3�������L���y���R�7�v�D+�is�ʹ3�{Ĺ�K���"�G_��6�:�9U�x3g�R,Q�.KI����
"%�d��2Y�Xm��pv�[@i�-�$m� 6=�����k�ZA�tز'��=L(��Ȏ��8ی��^Ko�*�}/U��m ��{���Gfɪ����b��K ��#�����/ԙ�8���"��>~��?zP%�<n!�[��<XT��3��i
kc��ݭ� �[�SM�bɳ$�>w��&
��=�(�z xf� |��=��=���y����0��k�JC2_ Ԑѳ����y���20�*��VA�6]
�С]ܻ}E��zh���Jpq��{d ?ƕ����8t��݄�r/Z˵�/���v|����a0a����Q%^����= �q\1e��F���䖑���۟d��2d^��r��6�S���G"��ӗw�F�݁1��gs��K��䛭�9\�� ����d԰=�i�f�,��msuލsʨ���P�>�;��t�d�?T�â�49��<2J��,YgϽ� �?��!��ZN�qG
'OJ�0
�{�E;��\|��M�OR��e�}]���Ln�m"OI�Ξ�((G�gk2���ٴ�g��x�-�_��L8^�r�>��x�Y<�H�D�.|$̭BG��"!��(DzUN�S�2�h~�:Ue�t�~����I�}K��.�����$$]�)Ɖ��PB�۞�(����n+vא�'qzJq�U���)O�)�Zٯ!��CvX�D���T���0���bP�g��eQ�'Og9E���tj�4Ý�f-{���X��y���yۥ��h��>��Gz@�΍B�ٻt��cO^0�"-<����r�.�����ဦ�̐�$8�ܙ4ojK�#Y26���]���~>����M�f._� fE�߷Uˇ�ah^k��[�T�i-�P=�.������iC�v�\��D�5����t`�r�Dƹ�]��s�����������0�k=�_�`�#C�������0�l���[�6�+U��e"��m�$�֣@(>�~9j
e����g�9߱|������`���2ш\3ɰ:�KS-4h<��U*/;���X%VW�YR����D�"iu�K6�)��7o��_�I��U/'crّ���q��{Ecz"���H��߿��﫺�Ǌz�E��	pX�U(b	{)Q�H@,ZyCn_hv�DD��M154*�8�MW���V@�:;0(9F�ʑ��p�����@���G	�<�kE�e�P�VI�\ڝ�a��)�}�A!	��i��ޚ�Y�衪�>����[u�7�潘���Ǎ�Iт�^�cd̠����MΑN]`V��?�Si����2�]�Рg/�N��"F�������������L�!���s�Vll=a1X��l��W�9}��ώem
M��A_m�,J_o�kV$B����i؂Ш�� t_��:�p��1;�J!G�'�̙��EO�`��"����P�ZR�b㭹���7A�ToΖ���|�\J32/�,��?�p�Eﳴ���nlm�k؋�ϥ�0��oi��A�5��]�Μ�����P0���g�ٰ݁�9�-M'�N_P����@~]i��Ԟ�������^��
1LvWQ���D.	�28]Y}�Ľ�6�@�b�>�bÐ.�1�_�W)�<�4�<��dà�xQ����C̭�z��+��&ԮO�.�ĝK*94;���%�wmOv;�Џ�1�P�}�R��x6U�����Gi�e��?��GG K6�mj% 3M��¥�<���%jC�����nQ�K����?Q��,8�Ǿ�Կ�n�a����$Kjt�?�����V��3=���Mڥ(�%�k��k�x�kT��`y}���'�:�s���A�����*XH���;8�;gv1���*z����*kU�[-U���<테h[LQ3��'Sd\8���Wn�Vgt{�<�\��o_K�W�Ͷ�!/}-��嫕�& ��2�5+����w�cFR�b�J�#͆1���}p�� ���A�;7����=��	0[�@���;��H���*�|�>���;
X�N��o˹Օ^��dDrt޼�I���9з��c}^:M!��fŌ]��fԤ9�Wo�	\)�ם�B��2<jz�4��aH��^��oP��i�@I}G��Ge��t��C����ԽP��)�ӐK�{�F��:`Z���f�(a~ݠ9���_��jc�׋t4<ETY�����	�1n��.d�s�@�Mr�u����r�W��d�rt���(f�$�PSx�q�B�wW[����g�uFZE��DOV[����N�)��b�b\�:2�Y���A^g�D���m�[d����1x(����=_`I�X�͟�����P��n�P-n�솉d
Y�r_a������o����{=Ȯ�"$4��� T�
�Y;��TN`.����񣤝c��zqT2��!; ��!#P{M4S��A-
��?_c����?+��4��1�U�dy�O����DJ�J�)��w�d����[���(�[g�Ho�����IN0[�>���q>�{�0�-�Fǒ��u>�N*���t���+��l ���@'���W/w$�����`�Z���b�iЍO��௮>��]
��&0��g�P={U(�ӀE��6-J�||"�6yCj�:���8\\!D�����T�>ZX�f�Č��hU�8�
-��'�*/��9�jq�U}�` b�6���8�`���;9x�̧d��&񦞧���{H���"c�2[i�>�I��<n�#
�l1��Q9�`e^PbKmhH�F��>5�2���E!&�,�5]�8���W���i��uX-��8�.e���t��9L�c#u�w�M��
��+�E��~(���bG� �+�D'�߮U�V�������/%$=1�nH�X���ME�i0�:�x���܏q2I1����Wq�-�# ��auL�2�#�j��[�����x�i(����ް<g��ۄ�şy��a�@ o�)�j����_P�.{�`����wĒ���c�-�K�>��3;�s�2a�yc�9c�㸥%��.	fS�yjyS�� �fd�8M{x�
��,tsݺ��#g�H����7���4D���i�q�Õ�$�7�cw1�GM
�Bj����MNs�o3�| {�������(z�9��/_�i�3�bjU>�#d�rw�fH�28��s��	��{�@�x�ӴD���O�68��R�ʊ�Г��P�E�Pٝ9��Ub ̈́Ht1�w`ھ����\%��mU�W������� u<S���C�Q]~���=��+�^�+Χ�\�t�t���[ps�иx��c��A�u�U�P��S�I���j}��!%���P�"�j�z�)A���^�^���INqs���	ѬY�1� �h}��N�l�U�~!Lj_��f�KJN�u@j��~hn��34_8S�^�*�����D�']���*:_���C��9��P��b��^-?��U�J�H��$L����'d��"�L�"A�`�����?V�9�a �;�2�R=�r�b�W�ڏ;l��X�1(�C��G�D���2�OoJ/@U�b��\�F�<���{���<���� M�Z��у�(H����5�g�n>K` �$2[+[[�L=M9�	�yy^�<4�$�ޕ��L�[7��lqI�⯹|��C�Uy��\&��˺��W�c�ػ`DQM����rˊ�X�]�qѼ��0�yz&����E��c`<��y�wQde%TZ������E8��Ċ��^�Ǩ�?����r�������,�!*�rhQ:N���]�0��Ǫj$����7��l��K�һb%��:KS�q�D6`�n1��.n��GF΅V��K#�>�8si������VR9�������v:U^j3�����[��Һ�6� �k<��)3W��Py�'B�8��>
��#=0w����� �%�e�K���3�I[=�h6ː�,8����+�2��~;�"��4D�5x���b��OjBh)�DViI�uP*X'Y�`��1\HtL�Gs��V�� i�ol�:B�����a
*
o���ݤ	'0Tm��p{�jo��7SN$y O�B�� Rc����o�A��lq�Bi�Gc��|� <����S�t��N8��9�T�0��w��db���	�J�z����? 8#yCwõ�Z	�r: *L��6X"�!rK�釔JX�I�
�<@�H�[�1��G-^p;c��O%��[���
|�ݻ��8���;�y�C�8|�R'Plk �W��.dǟ���������6;5�Ń9n(�ĞطV$dxq�ٞ�Kֈ��@^�/t������g{%	H?�Mr������|:T����v+��\��>̥C�����r��dȭc�l��t
.^����r��Jf������[�%M
H��8���4���Y���0+�D4��|��6�cc��VrHx.����G��Y���:)��M$�	��:'���@����o�|�����<��j�q�PZe��ȶ�H�Q�ٓ��F7�hND!b����3 =2�/f�Q��aRB�h^�R.P{<lm�Dy*T�Lj��X�"�(^����)�C��[����TG�Rq�ccD0��Ve�l�c�ϧR�v���E�A�C�������#�l�C0�?b��J��H��z����tY��w��`��B����>_|�^7o�����t4�p!�*��� X]D����s���ֶ0rAˎ�y���&�]l��]�'�,����c}1=�%a� K�E���R'w33ȫ�B�:�(�՜��=����9���ڻ=EY!0vQU�,���(\ء�G��@��
� ��/�U����!�AVS�����I�-֎��9�}�x
�e����r8鐘4��f�_�1*��)<V��2 �$g|�y��&q�bCP��)�&y�}R9�X���}KkC�v�$�-XQ��ԣT�	�脁��u��@����p���"�oe�dO�ә�_�ڀ�F�e!}z=�)�{�8�l{�*9�Fx���$�L�/��@���O�n5�d!��O S���`�J�;�#��3WKa�'7x�k%Rp�_�����)�L�	�vE� *:������"�9lfF��!]��׵��q{�ݾ"�H#PK7��#r,����T���(Z�;b2<ٶs�3(�P����2�!����F
��y�R�Y���T�#Hp�a�d[`lʇEX1B�3m� �+��U�͂'�5��҆�U�JZ��h���+�9^�Ĝj�%��yYR˞��&5�����(��_�>}��2�J�$�.$XM�I���c�j�\	��q|��i�s��gx���'�\J+�	�8��RX+��޺T�{2�t�O��|�g� I��F��Q3���I|l�g]��0E�b���p�	LT6$�B�8�0���qce/���	ֲ%xu�]`�]�W�Q�-Z�B#6�j	��?�|�3̧�F��I�I��@%�LTا�E�w��yrL^�@ƙ(q+��Wd�)�L��@N��������D��'=Zy�k7"���&'J����o!g���gr_�0�J���m$fh���Q����5\���>�Q�,�?V���GF���b*u
#�H�c/Iiab��de̲���N��_}��श4�dM� ?�����|�7��V(���D�|�-L!x/�]x6G�[m�;�>[1�L�j�q��3ppkZ8t��]U���0wdgO�<�0qO$��m����;��nX$>��CI̫:ۤ�?1����Du�Ic�9��оe�E¸d�����iI��(�����t38�d���}��C�xȜ�J����1����V�����z.��v�s����/4���6�Z���
�3b@c��3'��(�q�B��ۀ��k�9�Nɺz`X��کH�c7:~3��g=� ���4��}+����d����{����eCƞ�aw��LT��ud6��X��9Ӈ̣wq%����/��a�c0��Gr�%o�)�՛=m[]
-�����'qR;�z�]B!��\��K��qVZ�"0���vc�D=m5���%�'�9ss�H�<�z�EOK��I 6G��;�n|�OWWTp�΃9��#�\p�T�)?}Xs��_A�L�d �g�·���Q5C�)�9��ez�����#�8�ȵ�B�d�jҧh�fԛ�n�,��8���`�."q��c�
G7��7rw�x<�;��x�Z�1In��W½5�w7.?E1%�1���sC&�v슣T�<�%TE0����
������!�Ճ�fi�V%:�ʗ��ڬ��L��#K��"7W�� �77&]UMԧ&qt%Ov�����k�v��k�G���sr����O�Y��0{���i`[Hՠ<;&�9�yj��5!>�X =;V��؉����z�Ѫ�UqtD����'j,>�s���׫�=#"�W{#vr��'�qͬ�m��:MN�py��)�x�ј#j���1���G��(�h��'ݢ�hk��79;�먞����a�]�צAmQ�k,ϮU9[�E�i{���W�҇��Ux3�7�R���m])l���i��XiM����������TR�L�4ܳ����7�Thz�A�`��H,Z��h�bTJ��&�Y����w���aDߎw����j�=q�Ľ�����H�g�4˃��/� 3�e������@QH�#kF�u_4�C�ٟ�5u���	�#�W4A��"-+qPUF����K�n�i�P[$�p!�s�9����fR�a�,)߬V�s����tZ�q ;��8P��ɠ6HN�=G��TJ�I/���x��9I�fڢ���ӺE���!��E�x�!�q�K{r�Ѽ ��UUS5�p��!%b�#��osd4_刽�	zQ������s����]�]���c�8@|�X|��1(r��L��:��ESex7ӓ�B꜂j������m����E�F�.��L�xد��'vC/�,|��6B?c�����])�`Y`5�������v����<������~Lg�F���|�w�~;�r3I}���nҕ�((Ŗ��q�0�ܱ,4dZ�a^Q���z*�lFA$��W9]K��|ڃTy�,��v����X̮���7��#�Ƙ��eg�#�C����T�Yr~wT�?eͬB6��o��lP�j���z6CC�Vگ=-���2L�x�e*uX���o>��@ו ARL[�����$$�(������+	�z��>"D�W��5�f�ѭ ������XD�-n',AѾ*�N���N��$)�p�Md�'k�D�5�(��R�����%��8�]f����)`�)�㴋�P�\H���$�bV�+��l@z4�G�v�&͗:�����:��Ni6$��`.]�[�O@c��|ZPsHa@��u��}�����6ͨ曥*WsK��Z��(q�d���3�:��.@�qj��V�r��$�+�V��?�C=Hfڒ�#��l����kmT�k�gZcSY������U�9<��M��X��΂�h�uD��~$�3��0M��4�6�Z��+�E2��x���`q`�K
�Hw+N��Zč�Y[wN̵�y�e�'{�h���Y	PH@P/�j����0$�E�!Gm��IZ�qpĒ�/e�>�G=aި���yt:�seF�;e����F�eaj4�n=���!#K�a���+pl�}+�93t����)f���=~�g^�$�S�d�C%�}�v���1?g9h�yI1�NW���Ik�����p����0��)����dj��>�����8�%�U�fz���FV����B�z3��:�U<S�b04��
���DjCY��X����*���F�۝��^�j������?K`V&M���n��$�E��V7fP���Jx��>+�tU��u3˥�G�c����˭��,5��]K	��
�A��Ծ;%g�����c��]��{�9�P>\�����o 4�:s|���6]�u4ɌWT�4N�͵���uz�n·��i�hC�=6�����j�Mg�W�첊�K���P<����-�oe���a�iR�7�����;�J�W�X4YZO���"�݌�U�LBC�����@��o�sE_�xCc���301� �ee�*f��ۖO��&�K@��{�2�����׎0�ϸ� �����C�t�;3����MM7��v��0�
���n�]�^ޞ.e�G~v�*�	#�6��J���0߸Ɠg>w�e�7vw�9�PN�K(�p��+���Γ Q�:�,���S
������;�n.��J��MMn����Қ�m����g��)9}bH��BzqS����Cc'�}��6X��-q��z�~V�Z��E��\	�#zLS�b�;��OTBY�Ͱ�Ֆ9�
�$߉�$���/�.*\=�a�j
����q���<"�8��lK-&e>�]$���ʳ�2.���������e��3�o�ͦ�F��v��gt�D_�I`�r�)5(n%��2���qA�0�:���v���Ņ�*|�\k����5�g݇�`�F��n
N�RQ@���̉^EHg>^$^���ד6+��_���y
mc��>�<p�i
"��-��ɂ#��f'D�W�����-���S�Z`q5��N# ]us]f~�+8v/��Ҙ3	��yD�}
?hx���q20�?�wœ���dlߖԣv���Ԛ�^�荏�m%8Z+)q�Ky���A��$U-ܐ�-�F���=V��4��462�C{\4�� ��v���I�M�1��!jE>�I��_�4�B]��enp�*A�U�/!8��g�bu�%х[dy���B��#?_���IP����#ql[�Xv��gm��)�uGgF� �K��q;&w������>�;��fy�{n�G��ɀ��F��j�p�n�8E��As��oI�MR z�<�7]pt�����@m���u�O�aL���M*����0G.�1�N��w�RMߖA�� *��r�N���;���{~�i���2���jQފ���J�+�r�B$0]u�,1\��c�������`'�Q ?�O�4	�/�z	���`�gx����"<�A��Q�~/�S��F]o7���g��!k)iO)1G�To�=S�i�1ޡ"�H���>b~��`���N|�}4�{P�{��h�B>%��/\��5[I�s;���6ɽF:�t��re��͓�Mb�z~����F.ܟ��ۚ1R4S���`#�:PX�"u^&��߇�`J�c�8j5H��ٮ�MR�o��y,Zn+Ƙ��1���e�ȝ��R� �S%Ħ}���=$0<�<o�s�'N¾m����En��D�w��)i� �O?.�q�۟�E9��x"�,�Om�,Τ�����P�6X�qp�b��y�:c),;'�~H-�+���7K�ş��q�PS�T3�s^r].T�W4�4ƈw�_��w�Z%Bl(�VF-�R�yy�|K�]�UhSS��f<�&ي�ĝ���v	a�A?�:�*�`��S+�<1s�y���Ou'Ko�1���l��x��I�.�MF5���Ic5Ѣt�,���I�� G�D�v\|���#~���i�h���g�������u�Lw�`2^�� �����7�0N�q�h~�G�gHݡF�@S�u��S���p�1�gns+-���pa��|V�O5�>��7J��4;i62!��?�z��^��֚q�Q��0�%�r:�7�;H8���U�:��V8!�a�k�`ؼ��~t�&�C4�bwAE��m0$�a	X��dU=���p��d �p0P�� &` ���#<3Md���=;�$�	0�I�_j�[i��]��[�C���+���wK��a��<��<���T[��C����zĳ��8�[&��>m"����v�����6���Ac9���M��k�s�N���х@�w7�����qF��0��~ޅ.3u+�>w��̀�֜�`��N�Y��c���u�m�;��EH-���i���~ق5D�@y����Yđ�,#	n�.�1G	�Ta��L�V�G��JO�Jl��4T��j��7��k78�7��Y��!y
ΘÎ��
�\��Aɳp��9L�OL�|�k~[*u8\nxmg9s�Ԛ�g��h]X��NLG�&�}(P��=�IA?��uFPS�F�c�����-��}9�)%䨭�pȫpe�9,3e����9�|B(bk֔eǀ�<�mt��P����������� T����� ����=2h��.��}UJ���m��}�tL�k��4�{ _w�Nw���R���r�&�!eDA���ӌ����F8x*��i����bA=�BG�=�rCy�%?k��޼����Ւ�,p�5ݧ�:��`��p�ſ��s]��t���<���̌�����^qpq��l���8XӪeYm��D��@�����\U &�3�r�İ��R�7r.����m0�g��rj���&����ML��>a#5�$闯�?�Z��6V���c<�j�AM/	H�j}��۰��.l�B"�]5!�\_xh�f��;��5�U%��R��C�+��
���(�������m���E���*�g�m_�m݃�]�4I��NS���|s�QH�/V�2�<4��۟|�キ0�0�z�6�{ڏ\�_�����9�=��q�3_��D�bT��l�`Ύ/]�q��R撚:Ѻz�6�kEos��Vpfu5��Nݕ܎ߣr�"�莜��"�w���NNBrzE$
�!M��}�����"���nj_k�H ��~7[7	eu�{���	Z
Q�FZY�ԇ[�����L� �Ki��0�Ctݬ5����|�c�c�R�<�������z�}�4g�rt�s����;9�c��1*��yDmD0P��"�C�g��yE�+Ν����9(�3H+7}���~۠�q��&[�*�SiEG˞�7�B��Z�>}�ƨ����@nr<=Ļ�	��T/'�o����$�-���%V�V�:�8Oo�8Պ@���^�x K��ҩS��%���E�_o��|$И�r#o�Nï�a�<;EΪj�|e�"�w�l.�ˀ������T+"Y�=	�S�5�I�V-eg(S~ؐ�q�/��E�Oek�Fd�*���j�W�F�P��^m��bN�Ӳ¾��5��
��7�p��v5t7���6�A
)Z7u�{eq5��s��ej� u
�����݅%;�)1�)e��2l:��2fnA���!眰5��Jy(��+�K� %kޭ
�q��nU7�ϭ[ֲ ;Ʉ�n��K���<)�(��^8��tnQ����,\h; �)�����l����3�=fb�]?Ip�^��q-���0�����o���~1���8tvMD�[��矉g`��}��ޥ_�"�����r'x��!K������=�é���0�5�S�����F3����s�v��b�$�y���ˎ�W�:q�$R��elK�Y�i�v2�O��q'G��Q�b�}���9�w֕b���-���R1�pI�޾;��� ���$�&�#��`>�ٓdx�����eL�/�e�9ݗ�x{�h�6i�P&Wv_��b�LW�	�Rn��7
�|oA��ƚu������i@���pA
Q�,�ޭ����2߭�6��i�����r9��m���{Q͹����|�*G~ͱ���XsH@�Wa�4��˝>dlO>�d!�q�~��
}$������Z���-I/PF3�j�~`5�Q��{Ӟ2/�Bk�7W�(ꖓ}8/Z`�`�G��C��T�$5��┋�?)���W�T������L CR84z�ߖ�Իf#1�=�Qʏ��CBqy��|?V�f�.�^���<�V~@�&1�C��ٿTK�-L���3Ƞ% �n`?��ԫOs�E}��<��\,E�D@�Xm���N"J�y�e`�O:j
aEHц�n�5F�8G�P�}�
g�2���ي犿hX�y��WGq���j��S��?&S�+y��i�`>Ͱ6�~��uh���aQ3ാ��x�p�m�s����j�W��-j.��8�\)���Z/�࿑-��z-zXr��(fn��O�r��	߂�w�`ن���U��f'��ޣV�_z>�Kn�4�G�ӋdG�=+M��n��^q\g�aB���?�j�����x���-M�4@�=޸ǉϣ�^��!I~�%��N�џ[�9MQWc����vCk�$,���X�%d��5�����l5u!�s���<�ȷ�}w z�霕u��4��u07x����lfZ�R2.x�g]��T�Φ\�ݔ~GI�Զ���î���Z�Mu�מF8&����nu��V���mϽ��1���&�,��y�$�R䠳�4��qc8���j�5S�D�`�W����F�5}������6��ޜ8f��ߏX� � U%\�~�x��Zk;�z8�������CU��5������jT�d����� +���Y�l���V��Q�ا��B�4��aH��V�\g�>m���	2a���5�ۂ�O����R��) �A���s��l`�.N�����V*�㶖�bٕ���I�vB�k�?x����0R	��&Z��
��/��$0��@3�އ�{�0�[�Ə�����X����0$q(�2�4m&|�8ƫ\@�� #3��!T����̗�Q���2��KQBM(Ds���߿�D�1o��^�.�C|f�ɚ��D;��*j��+^��6w�{��!��
���ׄ��9v���Fc�1�LbR��A�M��݂zy��"�rqwb(�`�Ӑ��a��>����ߣ�:�� �$��~��K�;��5��;�s�|��["�1d�`=�a&"%����O��nmJ���T;��*�9�:mf���:�N�:85�p<�b�,>/�SPf�B'���>��+Xi藢��?��f�Xh>^$ػ}�q!|�9��1�E�%p�s­t������Ʀ�V`�@�Q_@� j\��Q�� kn�߽�/���(��E{���7P�?),�_B~C}�äv'�ac g�,�ʧ��"����Ϩ�#����M���h��q�#�(�p 8EP#Ʊ�!2	���W咥����c|\Z�h	�f�w|�W��,��w���Ni2������Xq�u./�b`FE�%Ԯ^�^
=�j#+��r�� ���\�ָڒ�%�TW~�>�(�ɹY�)`�e�)m�k�
c��V���iw���G�;�F�U�=Ɗ��W���5��Rt1d�')�� 9%2��� �C�}_�O���K�Ώ�4�˷���i�G�47n=��@��p�u-�㪭$hH���~^r��}�e^����B���n�7�G~L՞ڋ��+�v�&�7T��2�"�]����$�Qń]�>��R�@1������l�U��dk�(A��C'm0���^��@DE@�uZ &,I�>I,�J�洄�~ջѱ�њ��'����6os��+҇r�쨻�lǤ�.�h�so�H�t����S���K�m�&�S�� NB�l
є<���Bu� ����q�Dٺ��Iʕe���1�w}4���!��t�s\r~���z.p"n���%��3HǠ���wI��00�F�0�q�����hlp�z���k�ו�P�o��
�r�
�ۘEK�����P���(�:��`\��v��sVc*#��$��OԘ�SA�<�~z���L�Xҩ��y�+��8ŧ�q��>��O�*��*�qA���U˦|���F��};��|;��/ ��Q^��܏�U���Y�ԘJ��)1�L��K�&eҧ��ceƆu����!ޜ�az����6*���vE��<��|茶N��m��M �j�^f7��ס��2Rt][uK|�K9�,�m��L������XO��f%�q(^N����n�殩0w<zu�}��;Ê�0;)G�n�h�qo��b8cr���t�Tgq!�{�j�<�$!˫.	���c�ū�i��r�ٝ�7����G 'Iv�lrC�Y�c�(�e�}��R�7�ĪO\G���2حS%�~��nL�ϏF�����z��a�.JU�KE�����	�����q�42�Y����gO=��"�'�7$�̖�3����?KL݊*���$d���sѡ��3�:�Hj�K��Ԇ���B8�)�Pi��g�bkج��0�Z�Og�Z�'DZA���Q��9�������R�i�l�c�`g��d��+:W�H�O�'���Y��l�*�N��k�1bwۻ:g���1tӓ� wNIW�C�[��}_��?M8^5N0d�K���'�
����1/Y}��?!����R8�,�D�
	I�c�֍�D��R��]I�����9�P�8I�A��ܘq0����Ot���m�:����)5��Ȍ��u���ewy���@�Db ��п��D����BB�_f�tn���R��g�>�/��A�P�DAS�M>��(���_��׶uV��H
��Β�oZ����x���Ӈ\�xi��0'�ᙕg�~�5f؉4�� �B;�9��R�}CM��0ܷ"4ͳ>ý,�eK%��{���+_�@���WQT�Yy("�)@iȨ��X�Q	�P�����R��T��*�P��/��b�EK�� ��)7?1��G��F`o&F��g?ʷ���7��H��s3"R_f<��
�ˍ-���s� ��ʫ���[���3��*U@��F{x�,yp_
�)c�$� 6��#dG!�K�ˏ�,s�7g_�mKy�pi~�,�`��e|�89��Oڐ<? X��\�J�@��E��`^�;L�M��x�Ǫ1Ř�:-<�$ԔE�F���X���U����~�q�f��Z�!�mӍdA2�����E�I�����'9����#fŗ�,i��9*�ʘ$Q��;�s�reЄ9;A��|��e�AS_��GkR1��:3}&o��_��Қ��iVU�7�~�V2��MAk�����/9�?!Ih�3���yx#�+����*�|u�c,�d(ؑ 9k�id�/��7&��T0��H�!�YG�rz�E���0���=*x,�"?��ԙA6�h'Hv̹ƒ]q'�Ѽ����c}N�S���Gi]S��p�Q�B�]6O��]��t��K�o�!_f��emkA�s���/Y�'�L��y�0�F��G��A䓖�ʴ�s^�@�����F�U �d���J@8�ډ�8�]��K6iLH0H��s@��N�Z�1w�೷u���>^�Q�Q�2�����,��v�!�)�o��R�(dhhF���b��L�.�f�pٺ4���_��
�����*���c,��ѓ�ZA)�� �BO2��%	���q�4�{	a]M� Ef�%��I^@]���k������rFԪ�ZW81���y�y]W��#��?�-W��4���5�{9���0jm,;�����O��X�V�J�l<��<���!|��r�e��A3[��%�z��B��fX 	�-ˀ�/��k��M�	���.���V�<\�9%V$*�IWAٝ���ֽi�ߩ�<؀'d`J����G���%�pP'�����e�\ao���=�Z>�>��x�۩���rb��,|��Y��'P��-u4�|�/_h��4;M������$����L/�%}�A��V�%���~�
e�M�ADs�ךu�,� � �r9v�Q8f�j�r^c��~����$P��n./�V�W��kE�x*f����Z�u�R�����Ί,�FQR`)`�-��O�U���s����I��w�N"SX�o�����}(����@]��U�u0_�.�.�"�N���Y��EUZ��@��1��"��F�M���?5��0ދ��Y=%�U�[�1\���
��1a�����:�P���+�=^�)�硣HM�93h��!	�C�����}��,l���9��%��T儰���o��$�TWR�n���GюÔ�ܺv��3�7�^����[��|�܃C�4��h����ȧ����	�L���	��ށ��*�ӟ�)ۃ��9�#��=J�M*s�+*MqX` ��$�u;o,B�\7ӒP<7�Rd�h�+5�
`�>G~\��l��/r��,rJ���b]�.�o������1���l���ҞD�3��$��!� ��GJf������)tw'@�0t�:�#��͘���D�C|Q���ر������S��Lg�o��b�B�G�*lp��Lv�����F#~b]�#߽����X�*˅���� V�>��:}qp�,N�7i3;'4i~&I���X������(����h��k���A���-@�X|�"h�+��]���|g�Aw6�=��L��-s[�����JT�^�Ґ�Z
��t�8!�Q�|���e΋W$��b�p����N"��`}������*��C�#�4e���W���K Zƺ��8!(E�*g����}��-�	�
K$o��CP�d����c�^w��j�йU���-�3;D8���TQb�҆1_W鲹Y�2|X*.zf�$�ږ
�X�nJ7�O13��r� d�%wp�np�������hLc{5����P�{��V�q�%�۹���&
u��˟��hf\"*�g���*��RQ�i�h!��C��l���ެ���'���=D��C֍�[R��t�s�`���ϰ&sA�;OE[���n3���E�����r��PC!�2����]<��fa�;�L3Im�~��y�)��5����2mq
S�/�2G�����x!T�����8)�pT�O]��>�z����jT��:��y{���i�=�����򺷇��ƣ���Z�Xx��%���]����h��=���v�Z�G��q?�L��$#ϞvC�\1���}�{P��y=�i�����+�,��'����3���U|���+R�l�jh�!Qޕ�[c�H�=Y{x�E�ϣczx�[�{�k�'Ai�U����-.�2�yn����7� ��It�z=K�){��εAoXb)���a�~�v�@�B���H�� ���6�4�{d恩�������aiu4���G�t�'[�A��t���чBB~��q�-��/9�������o�ý���qÌ�����v����Ȳ'�����p|Drr���	�J�ڍ.�)�8��E\�/���/z�2�US�˾���Vw5�_�E��i���޶ �4U)��n�^��9]��|�7�b�I\�R���lsB����Fr �FO�� ���ֻ�L�#)#��a������I���,�mr���J>d�����ѻ��a2;�M�rj�{�g�AVO�L��x���F�~�ʽUL&�Z�SK;PcUB��,q��c�N�0�{��G�>?����6Gb��˺�I	�I|�L�Ƕ��ܔ<������,����h6>��a���1t��ڸ@P�؛K�Θ���u4�EA6���Y��"���;;����'KK���� 7m�%�_��v��0�8���"M�� ���ǹr���f�t�L�:�P�gS�a+<ъ�z޹�-�`i!-�BT�B�i�y�r���p�/iIz
���^�Ϣ�e�g�ʡ~�r�kVHD�*���MC�� �L�Z`�ұ]9�0ɜ[�%��(���J�<=K�[N���8�C��o�D�I��xK-�s��*����{���$�D��ar�3]��˻G�=D%��몃2k<5��cﮪƨMѪ�&�f�Q�A�ERN�T.,��oUWzL�Ey}4��`*�T�t�{Q�d�[�5�tsTi���!���A�B��%�?)��L�~a�TH
{�I���Eev�W��Z�8�_�4b6HF��\�ϑ��_�\�
m�Oj��}��pŬ�fu�X�W��S�
;�b^�ݛ8�W)���e!�=�9������$���sYT� >=�j����m
F-ߔf�raV���%������,{�ע��v���V~����2�*�h�Rs�E����w��<J[.P���1�I�DI��r]=�Ẽ�9F)��9H�rʂ:ѡ�)*"p��T�H�~����o}�ԾQ7�4Is��ʦ<�b>�`�u����Ѵ�?�G+)ۮ�L�k}2�GW��8��9@!��1/�sR(5|G4�������X�D?�r�E_>6x.SK�p���{csԀ��#�5q�һ���ffmc%��^�-d�����ɋ8���f�M��	W�ⶭq�<���+��0��I%D�%2I���D���8}���p�:k �`}w��~\]�J�Jt$��ǟ(�Gg;e���c�f�my��Öp_��$ҟ����KT�y�U_Z��Ʋ��=dD6����+��+�I76F�@���3b�L�EYB�V~�> D%IJ��]ȋH����)�� ����(�����R��m���>$���$��63����'����v��'C�їMH�� �
Hc��o�_Q�z��ܳ+�C�c��49�7R�٥%�{�P T�����*�����HS�G�;Z�ljC����_���C]��T�b���=m�m���%oHY�H'���PA�������v'�y�Ǹټ�蔆�j	�B�(3;u�^�Ql��0$���5$��&��G1�J�����d�
�n&�r3x=z��U�h��>}:'� ��fCFֶ������*AQ��$�|cނK�r���BRVNS�����@�E4����Ҍ.B��2�1�$VL�*�?f_g?'z�$��ZՌ��L��InkI��m��_�7o[pT����T�q'�4�~� s�SԪDo��Q����\\������6΢���Pm�����Z�����8:y�+��0��Z�S�΍���[pl�v)HDrb�L8�4�>ĺ�`,�M�@����'�W7/_a�eC��Ҫ���͗��}��h�`�Sހ%�[|ֽ�!�-ʹ��A5Y�}�N��!��XB��J��gq����$�����S�(��ש>@�0�JeU�N�]K���ߏ��>�m���_��Χ
��'2{���N�
��D�e�^Y&)���b�����x��%�w�%�����Ce׋��Y1�"yl����c�%�O�9��}��}IH�5J;��EYC�.m2�Q��e�����4���I��˼hi#��z��~�1�-5��5Pɚ5���Z�2C�e>tJP�a!e��W�}e�I��i��F��ǚ��|�-xG�ݍm�ئwK?���k�Ea}p�Y0�=�	��;K�x��^�5��O�T�I�l�F9�?�L�Jb�Y?���f`̧jI�����q�O�e)�@�8�:�8�ʓ$�7Fv� j�e+�{p�'iS�XS>}�o�61`����3~#1�0�&�q]��ƑSǵ��'�r)c�.ċ���L&|�|w�rV~ya��o�U�Q�{}8�_�'�-��S���0&��Ȗ�7�;g�J
,\�3��EO�����0Y�"$�Ms��� ���x0A�-��]]��rG��(/�8UI�hP�.�d[�F0�$���Ҹjw� �A?n�fm#�o
8H�$�8[�!V�!���f����/m���x��A���|^4c�;]���sO�^ �C�NM�]ʽ�ci��As�&Tt�'*p!�I����J#��A��g:����t�友�%;�B-����-����e^�ц�W<��n�DYњ�X�1������]ZC�5��?&�_pN��[2Mć�X�EƷ��@o��;,�	_�����zs�؏㞊Y��w;g7���T;f��]�cZɵރհ���.�/њ�ϊ�y{�����^Y �ǹu#
 �����^Z��?�;���U�U��i��i���^g� o�=�
lw�	y7^�h#A'��,���fY��'BeLB�'>,�^$�
�P�޺J(��{U�D�:�Y�$r�N)4�7U�'�]���[𼯴Ђ��!��.0ws�u�����	%�I���3���PN��u��x�5�^��͊��I���N�z�>����}	���X���;�*٢Z��?���X�]��'>�_g6��,l���F�$�=�W�zb���]��Ż���׼$=t/�ki�����﮹�������Q'%
6������a�E�Lx�	}�����A;��C!g~�$�uH��9��]8��{
�@U9����g�ݴje�A
�z�1��_5|�mb����~+�[5������s�P�$4^ﶶ~���{�ߧM�]�I���k:�ӆ\�x�56Nq	;2��&���.SV�-�|;۟��E�\��,3.X\�M�R�����9��P_�bXrd;�����G#�#լ�Y���O����Ql��"�ܯǪ�<�ףZ���"��n�	
�3�}���*x�y��`5ɔ�$��z��@0X�Kڭ3����<��Y���B	&4P��aJ��!T�Z��^�!ۼ)����\� ����c���<�J��� ��x����i�|���}�Ґ5w�TC]؜=�j��p�� IkI�����g!�?�$tK��t��%i1+�S$_�`+�F��Mߢ���o�����ISx�׊��(�yY$�b��A�%��?L�TW�ks���D�%|rz^(����x�9V+(�8S�c��F�C�	a�e��%�ܶ�6mC�^]�+�|k"y��pF�Ad���n"��,4Ȏ,^A(zu�Ax ��`
�~NA���&e=��c�HAv�B�B�����ʹ�4�� ��7� 4����z���t��	����%H���Y޴Qé��jx�}���u������x1�8E�1�z
�����@�~�ˀd�D�fM��ou��I\D��fN*�Xq={*b�٩洳�<�C�Q���3�~,��9�������q${9A����a+׉=0���.��1lKk��,Qe�K��r)��du�`4��E��<_��{ڇt_�e�JKĀ����C:`����o� ��f؉d� ��9cI���=�|6����ޚcX]�H�݁Z�'5�n����{�0�d�oh`�+﬈����4p�D����E�A���b2��vȢi%�;'�Mh��lޚ�hfd���>�P��0z���u%EI��#�,0��B;��#���s����m�'���Eқ��v�KY��솣��[V��?B(-��"dj��Xem �	�M���#b��W��(u��-#J��.V4�>)�����ȿfWT[��ε`0��Ds6���!��2h� Qy5= "�#�w���.	Uu�@۟E^F?&�DV/De����$ Bw¸�M,���R�e�W�b'ʱ� ��Q�z����Y���2Π��YI,�\^_��R�_�uik]�t��@����Yw�3��I��9ҫ�	�ӱ�q�9�P#�������� �I$nr�cI��Ť !F��#U��;����E��i{�����K��N7�H8u�X�p?#ӡ�W}6�Z�k 7!��t�����ܙu*�ښTH�Ȯ6���?���+����h��a��&��-K"��Pw����"���;��i��I؇�DoW�m�_��ޅ�	�2��4�n��	���'�Y�4��6'�Lta�kC������1�z�5M|�G�q\X���_���юm˓l����l���K;D|�g�8,�-���o{�@��k�;����ߌR݉��C�!����48l�����'����>�cH[�ds�y�5�����N�G���HV\��:����9�f ��!pG���0�E�����P螎s�;Kw������_v\�6k����@��T��Q�\���՚@��I����ZH�@b��Z�:�����<>l�vA���6�@�q�-1v�O�	��֍[��ޮR�[Q�O����唞M�� ��~4�<(t()����C���iJ��>���n�r�
���8���}�Y<���W�xT�DM�V���|�5���CV8��@�Գ�y-4ЇE0qݮ�.넮hi�|�|�'���	]P�e2s]��~`FA	�͞�wٌ�i�y_2{�p��9 �No�*�JS�P���)���U�[����XM�&�p����?+��2��eI�:`�S���X>�~���n}%~ò��pFj���j�LM���:�/����Z~����N����K:���D7m�p��{�^�O�l�3bE*=]��Pf�����Ov:`/��q)�*j�q��[e�g�H���9;�1�!3]c������7R��N0U=�u��޽=�0'e�;���e��������?�k��5j���'A�����{��9� ɪ���a6��(z��1P�,��uo�\t^R�^(��e�)��U��y:ezy�+�n��rHn�~`����®����6<c;��q���|h��*���vc�a�mQ�ٮ� I����XЖ�Y�g)���j��o|1<8*X(�ZHb�yi���|71���b)ŪHr/u,=�(r'X�o~?�Q[�=��_�����-�W�a�:9��汲��I�e0�^��^x������x�ܬ��
sP<����T�Z�xN6Oe�/���^w�d�nl|^V�Wl��8V;�-��W�m|f}��$� ����N�4ʑ������@P</�Y�O�o}�Q^S��2��v
:/T: �����Q�[�'y{�v岝�#��o���m��,�]ڐ��J�a���p���̬��Bٵ�U���RU�B�'���z�|1���	KG&�8A�^��Պ���W'ƞ�?ze�w�q����_��ׄ*��.8GߐA������8����R�z^/|��8X
N��[� �s97�\𤅲.6_b�%!J'�;&?i 
k�G�Qm���ǧ0޾����T7�w��z���=��j��i�N�v���/���M� :ȿ��VJュ�You�h#�<���]��Oŏ�m͊B��sO���M�0���� ���J�_�>[A��}J�p��m�bK7�>~x�ޕ@5#�|�RDf�x�(XS:���b#�w�;⇬�K��A��z���?:.q'�ƞ�^mP�z@�,I���"U�XI��(��A�I-��l	 ޝ�r��5W�r%���e|�����]��`�E{��	Hj/	H��+n�h@��$N"Ђ����[[D�ܫC�[C��W��|z�f<��]9a;�i��w�Oʏ
�σ��7��y�n�Gܲ�jؠ/0%�.|���"gU��;�Ì�[C)S�2��Hk��hɸq��8����%LqІ��M�L1�����ݞ��8�
�\����KJ��'h�A��w���C�6���Y0*RB��i�U���=�Ǭ�*q[%8iS�}s�vdz�u�[� �O��
�t�s�Q�m_:!Ҳ���2�>���Xt��H� v{�4{Y�K��x����_"��Z�t�@�ʜ��� Id��1��H�`����5U��yR������0���\�[�g7҉��}sr%�d����?�����0�s��z��Wq'~����'���vЀ;*��,���h�.B�Mm��x8��O)74��R�BM1�ק���b��$���=f��M���gkljN���MK��tD%�<��0B��X�����	��D���򫚆 �B/�Jfז(�n��꿺��OK�rt媷�� �Eʤv8t�2N�7�򫂽@/��\Ȫ���x[����1=~^�K�!���Ia-� ��&�P$�d����8
�$�k��� Z�l���O,��h@eɠZ9bY�w����ϑ\�,�6�T�O������;}���!|��@�q�ųTti�뭎-9�N�L]�(�=r���M����G0⿠�3݁9�>5m
Y�ۙ�>�h%�a�ݡ~p�F<+٘�,rRH����]X���]'�c���>R�Z�,7�\�I���_W{�|�V{ ���b��ch�����R\ݾ�NJDAn�n���'����⨫����M�-&�f����eO�T������8�Q�rD��/I�T�I7� k(��L��"6|�C���*˥D��z��|�٤[�`s��rٶ�h�Pq���׬d�9hw�bu�659��G�����̜��i[���
���
��R���qn39]F��h�_B�a���/��|H�Y�Cq�_(����� j�p�1yb��o�O^~�!3gXB�D��4��X�p���8����iB:��Y|؟&{pG"64W��,�YV4Z�`R/{!Ms��	,�h�V
k���LRq�w�[bB4����z�.��ݱA�F��	��8A������1�k��p�O�+I,H��X�pE0x��i���C��[����iᴋ.�6U��g�_m�_3��Vwz���Q
�Յ�߾عőf^6a{����6�Q��i�zK�����n��Q쯪����+~�S���g���ݢ���#�Z(������EE
/b.~�9)��,����'���PG�3����!���YBF�o2�-gH?S0�Dt;�c(PJЧǁ�mk8��� �XN�Y�R��+��0_Y���̓�BM�:��ٔxp��t��*�<B�{M��>��q�qK�2]��]���q~�C]s��}�)=6s�p�g��wX�y\L]�O�L��\�N�����yؤ����C�j��m�?`��Ϫ:V��^�	�����FD�<�]�/ɍD�}�+�	l��;w\�7�ۛrIJ���c#�&�%$0�manE��,�H���D�A.�4s�O�u �>�7nWo��G{�6�/�]��ƀ@\枹���.��i�� �0��G�)�u%2"�f!W6�-(;�'�]���!��)I�$���kN��R� l��R�4�($�8d���݈v�z
s�'�jhtz��	s�0[����c��xWĢ���P���#����?8'�&��2*R�zޅ��ԋ�����ԛ���l�m���o\�K�r�6��u��׹�bYA��~�A�\���'Q������P=ԭ�22��DxԐ�0��F�s��;ndx��t�15X�,�����$W��hK:R���P2I��X-[;�+۩k����(����~p���y��yi�Q�R1��N3���l'Y3�,.VBX�'2����11�a���٠���_�����<���c?N�����M%�}��gs��b��h:&�F�t�����m松M�0�`��\��|��g���
����_l�}��@16�l�������4!?�WmNɻ�9l��^��3]˺���|e�n��'-PW�Μ�f=�a��0[��]�b��۶������3����d9:����]��(��=�82�jf�qz;*�<�y=^���W��G�|�Xoɾ3�ף�PYP�s����똖�1i�+V�q�]3�;�rWM���蠘���B꤬��5�M|��t@��$̰�����O��P=��"�X��e�{vI�(���|X ��p���֐p�D��ib{�ۏ��5�ٲbIk��tIխ=�o��>�Y�A�a�{Iى�^V	�B���Q�P����m�GC������6�u�8�H�^쇡��ʛp�]r��nU��]ϝ�h}�݉�2�uvsG���>աx� h�������!D���+:��u��T�`��g�3��q���ٱO��}��2�L��n)V�]�-�!"�X��t&�M?��c�����α�e
�d�,�P�s�T�1k�����ƃ0��='L5�ƜϪ��=�,���f<Q/�_!i٩�.m"<7�p��D>��n�͂� ��~����:���5���ֿ��Z6F�I*�ۇ�9K��bt��a�kD���D���*3���-MiR�ZR䚬��E�]���W���	��~y��	ҍ���`��'���'
:��Q�\ӊzEE���)���Ȟ&�E��A�0B��6v����-�^�+K�!�k9�Kg�MzO���g��=&f}]�F�Al�,�gg5'm�l"c���*�������Q"��9�p~D�v�@��l����r�^��/�I���H���S���p�
����F�r�^�T${��]͉��(����P&��N���"	J�4�'n�w؍����@��ס߸�5ZRt�m�k�ٞ���wb�Ҳ_6���KĜ{b����¯^���B���h�a��O%0���U��_:�>C:�ٷ����F	U�z�*-�U���c"J0����ƐjԵ܉�k7^Y��qzq�N��1�L!.��|��չ��7�D{�AY�����5�F�5!��3�T����[����zp�k~�)���+�l�u�#�b�^�b� ���3��O��0D�u׭�f���L9}���=��
�W�bp���E�!�\���8Ǣ&�	m�
�|ʩ,ۺت�e?q��S;����7�gtD!��I�%-�Z��W���fv��5|���Sep=ۺ'B}^O1Ƿ�$f��<z}BG�y	1�LǠ߄!���]hO�Є�z����s,��s�1�bM5�bٱ����ˆ5w��<c����Uc��.GpO8ş=H� {V�<-},G�o'D���q'���UR˒�_�͚�W$�E���,��y�g��,�C3�g�S'�
։u�P�k!ǯ��/�c�G��S@.��@����9W�O�����w������/�y�,nmRe]�jl����h���9�����+Ǡ��ЗA����[Z̙�Ie5��dEML��
0�leO�c��,��Ӗ�f?�M��*8|�U֢ 3~ɣ��VjLu旺���d����ѹ����J���а&��?�� |> �͖U	�6,�]u~{=�����!6�(�"	\/�Q5�6LDf����M=B��w����=�����o  ��H�����6�;�`z��s�Y����������P
���m\A�x��Oaʊ*�3��F)?� hk�����K�,$e-p�@��Y\s݃�׸��jW��IoA���Z��PA��bE�k����5�b���q�K�l�S'�I�U���F��9rE��
��M�m��5n�L�ck��wߐ�hӇ��[����C���
���L��E�Cs���Q�X�L���:��e�Xڥ��`�����5v�K�����u��d�*A���Ѱ]����9�G+I�?�cͪCҠ[-��"�j�T�~Ƀ��H4���iڹKrtX5�%y��g�~\��,�c]�;譶�~�C@M��Q=1$��32��lkI�#"��?���:��Oص���R�Hl��?�6ݍ��N��i��{d�Nd=�"�h�`hYX�����5��'?�c{��9�@���D;�A�rQڈ�+s���6Du����LpN䗥Y�+��-�lH�H�j�4����Wr4��Q��lx_�u�5�z����^	�(7pZ��5���ݚ��2��7_@�����Jh=F��@kx�0Y�7�Y�p�����kAԔ@��U?b�"���O{�7y���ew�\y��^]�������wj�(��y"u����ߩ,3�@���!߂r�#�EĻO�^`>�yb>����Zg9�P	�^���@j����ys���	�g]1��35Lu	t(����赳�/�������+�ܚ� ��n�4�ԭ�G���Ԧ;U���JA���e�q�)����<�'g��h�5G��t-$$�e�r^��_�MT��'hvY1��F"�����Q�XT.��ݶ)0�)ܖ�V,���|��H12����o)�a��)�+I���W[�3$�t�tcpd���/�՚�9A�p��0����J���1NQ��%���,�u�Ӊw��+��x�]� 8�5R�	3=������RB4�TM5tU*�K ��M��� Qy�%�˖��dy�$�p�D��s���Ҙ��!���.�_�0l�g���#��P�ND�Sb4����^�xD���ץ9�%'\��(��K��#W�[+!���V`����h�3���O<��b�����R�����C&N;�&�ጃSjSB #c˙�QF��(��#��D�.%��F`1�U�Qp�y'
�C]�y�z�I�B�dZ���,�m�ؤ�=�����$���C��Z��_8GS{����c�R��	0A�]�,=�WcXo�,ͷq�h��ͫ�x�K��B�EI5�Z�����?�h��S
�Sbg�7\�z735��Z�K�����H"���͵i,�׋Ҧ�G��3F�NʚG�f�I\�zuZ��논�懤��&�i�Z(8W�<��?���<�s4%$U��0cB��6����t�X�|�Y��E� ��{�2ڄ��aۃː���8��������N�9?�|֞�ot��ਯ��u���L�Mn�rO��|�K���ݾ��w��{vug�	�0�?�>�`��m7��:D��( �ք�zl�%7%�������T���xCk7��[�u��?�$�&G+�O�}qf:c�!�9V�)�H?f�!͠�I�?Ω=l�?�����*�%f"K;~�Ԏ�ꮚ�6ѣ�bÃ��_w���~�y�V�;R��'�'��ℋ��f��&���_"a�o�F��(����gc��0�ɀ�N�C,{w L�r�ʅ~�HW4O���։l�]� �Yo;���`bף�TjH-��_ޡ7���M\��6_X&[�$%�g�dk�$�R�dA�V���8�-#Y�:ag |A�C:p���Lb�5~��-�o�	�ܭ��ʨJqc��q�ϲs�p`A�"�o�NAᩅ@�(����� ��L�w5Y>]��y�e��F^$��5-��f�Z��+^�2~V�}K���i��N`d�w9#��L(�Qx��*0�Ŋ����|�H�2�)�%�+<��eFUp�����>,��c�h��g� ���M� Yk��q�bL姗������Ҙ^`�9�u2�0.ɗ��|#z�<$�uY#���ƙ�sn)��ͭ��
��i%�����ب��3Lo�N.H­��d�5�k\Kd���8�`80Rn�Q��ؔ�$c�iބu�w���	����e����^�9��=�����bu@���!2|U��Q�2������?kơᱱP�K�KB���2�6*�,� ťJj�X}%,�p0�Ք^_p3��KpWm��L/J	d:`�`����@܃���U2���^��ݼw�f+�VV:>+j;gx�H�!���1�hh�K,���0S�0��5�%��On�C�)6�f��.5z��+�"y�2A�;P�Ez�W\k���e������F'	�@!��3��
��6\�^h�o��G����{WXT��nPĸ���z����#��=�	�@�a�� N�GI�G�di�A&�V��IM8ñc�FP�-33��!�4�N8[J���a�����I��Ӆ섨�P
&ZMQ���^*�`��~����7]�Ƅ*�͵����||<�r�f ��c�f�o�Oi�Z�z�{,hU�OQ͋�Z�{�b�+�v��s:!G����9i��iukF]y��(ɒP
��5�A��7�8G>��Z�S���p���HQn-/�g�-����Q��3J�G�6]B葿��_�*ְOs�D缭%���=a_��
 ~,�	M�WvȪ80Z�+���KĿv;�j�	��%��������j��<<���֊P��A���+9h�_���~�_%��MǍ	�oHc�|���5�b?[�̓�"��o��f��r��B��㈤G��!�n�����2�kٱ��~�5T��<H*ih�я<�u�&����С�WR#�ö�;�(��g�)$��H Ah��aZo���X���)Gk��̡��z��nxۃ�vP���B�$֌��0]�!�iІ����m㮦&��;���jն�����(��x:#��_�o]��1�N[�&��o@��K�=� -A4,�cN�.�{"y��A�R����g�B�Bk�0�����F|�$2ZPXMf�M��ďq"�x����k�g�"��6����NQ���rD(ijN���,�f)G�<�7+���M"�dn5��YHT�������?������0�Ql97�JF��ܰ]�5�nps���d�*N����Gn(���|��q�mbY����^����]O�+�g��M�Km�����<�YZF�a}nx�\8]���JW��ql)�e����?���!�h[��{��p�x���"X�f��I�1�mu�]3��I`�B��A��p��81��LL�\{����ņzQm5�#���Q	�+0=���r4gҋ�J��ʳ��􊕲t�bJFܪ���s�x\�	�%���2^�P:�ل��!!���A��;i�`X�oTԥx�:���_$�kM�D�:�ώG�hQ��2���Q؇PW�n�ɖR�<���SŘ�h��[���@�F'��Q��-�х/*��·~�B/�ś�+N��C�����Qr��{�:��j���Y���!�׵4��,�t�C�����)�&��
�/��������R?{�YC���|��JaC�����ݿ
�#�m�IQ�J2�����o���i�jp�J������W��-�S���:ﲨa~�'<���@�#��V�X�Y��p�j��A���c�xNHѭo��"{UM����
r��7�d��2b֨�Q�ƈ�~�0�|�ަ�u6��R����h��j=����J_ZM���=\&���/���-���$��Z���������_S���W{���x��%NL�F��bV���(�wԦ2��P��v����th�@�2�2.l}\�'i�G�:��@����g m�:ZܕJ���fΗf>[�b
 �$�|��m��} �O����dݐ�a�g�j����V��R%ԅ!�?zF�wO�M���j���K#���Sx���8ü/X�ܽN�5��ʈ4֌Ec�do�c*�jZ-����U�2׾~���I�{�GnS�ug��O��EO�XDm�@_F����d��L��D��M�f?�]������o$�e��,��xO��t�T�˻j�*�$�	��=�C)?
n��!�xvצ �2E*�v��v� �d-���8lCQ�����l_���/����sCI [=V�����E�7U�:�`1�`Ueg_%v�zS�2�����%1�;����
$����*�n�(�ѭ�y�1 � ��j��}�<��[�0.�p�mU��e� f%+�h+�����f|�[J�������c�68P9ӛ�wg�d��3G�Z�>�7�E2D����*��I��䍲�@� �_���f�����G�,E�-�L� ��'�H���3Zl+��J���Z�i��Kg���-�3&ó� ��k�0 ���K[D@l(t��~g�h��&�YZ����:B�B���~(i�o7U��]�4��rFD���'G�E.ҧ�\6�D\��x��'���X]L�4�-X�7�E��v�V.ε�d"���y��q����F~�DXS4�!@fԔ�g(r]�U��0��Q���'ˏ(|����Z������,�� edp?�)t�dS�`��N���?�Lu��0\��9��~Ԅ3�d&�m�De^!����
�(��i����1ߜ�����T�Ea�(��kH��2�k;�f�Ĭ}�7�1��d�ʉ`�I8{�=�4����7]����"�գ�}���tC!/�%$�Qs�W(��2����k�۱ڸ���<���Ɵ�9�&�ra�KP>��}�k�o~X#_���9Y�������z��ݬ:e��[�.G�Y�� �^�Rqs�9]������iND��d /9���X
&�^�@��=ks�Dp��L�W�\�[�LB�y�wu��S�>UJ|h������r2����LJ�Ii�<�l�6� ql��uW51B�C�HVj�����_�^I�(����b�2���S�֤n=��"�b�Ln؛3�dM�*���~s��Ey�*k2	�cs�
`j�Gr�n#-
�1��{	�G`�h%������~�E>%D�3���y�7��-�Ϋ�,$�2|�,}#�]�r9?p$݉l7#N�;���*"���6�K#ڟ��5�6*�c%U��xep;��|�))����^H��Dr����+=�@�z�E���w,o�J����5 �[���ӎ�λ�-	0^Fȿ
��L�11{�~�F6$w��O��J.5o�oA��w��z C�w�d�O�:M�!ք%}Ww�����+,�N���B����|h�Z���^��w#���پ	�0�s���EF-���h8j���Ӡ���&��i ����Ð����=o���B��Un��d[���'���N���'�B����N�;@���=�+d��L���F��d,�kmH�~j��u��g<���&�A��"� Ք,�A@:��֔b�%v����lC�F��Ⱦ��D�}f��\4ŏ�
�B����o��[�F@�]9��:�XJ��[��s����+ng�حq�6Y���m��.��Y�=Ā���^T�O:*x�A�%Q�/m�[~M�z^z�E�ñFR���e�\W���_�$P<�����������tS=^D�f����ch	c�H%L��q���Pg]���ϩ�dW��i�#ޔ�Я��
�\B�U���m�9��ؗa_$�{6�v)V��a� ����l���[�ѥ�y)���EB��1[�V�<B�*�>n��1m nؤY��,�a4$p�!b�G�>0�o�	�Q��_����]�L-|��Jo�.�~�^�ʷQ������bR7i*��B ���_��{�07x7�.��M�r���l�
�1���s=K�R�\�׾�E�2"��8���_W�D�[��C���i6�t����U] ^������'�� 7�e�����k�קϤ�?j�zL"}V/k�P?����r�aG#h�h��Ǧ4x���#�Ls�c��74�-��~����b��6`�ى����V�d>g,���̤�Ė�U��C(	�%�2�^�M�8��������+ɞ��Z�t��/�s��q'��ӷ�޳.Uc��E��dc��\��㹬�d��xR����fwѓ�( +$SM�P#����9h�df;��Ѳq�����1p�z����u��iC�bg7ɬ���� �����{�6���_�az�O������5��Z���*�-�i5��XwZ�L?�0�z�C������hYzU���`��Ġ[K%��?~ma"��ACl�Q�4H��D�}êI�Y27�����N|�m �̀_�eЗj���Ù+������ƦG��������XE�sZ�Vl���� �^��~�!�ij#ɤA󝝇�l�<̈��K�I�>V,����Q%jo����Z.n|��ԧ�J��
���]&����TFo���'�GxQd��M"c.��4��������׹l|kO�R�6<�2�����P_�d��0S�0���w�+�� "m#��B��+�R�}�/Yd����|�((����NZJ��*{������S�o7�,6��A�$,����9^�]c��lX�+˟$i�Υ{��;6!��B�v�!꣙�m+mT�x�o�	Z���$����-��rAEu�{�($X�������뭶��n2�n�؏}b�eVa���p����`}E|"Εi���-�����Q:�'xZ��~[�ʄx>4�����!ϑ~�^�;Wg�Q7��f��6
�X�ݗ�g�q$�	]~��@�B��t�r���%�ZG���Yw�lI�+7D��t�u�֮���:6�|v�����c�!U�Q�	��h������<���`'9Kg��������X�M�����c�@��J&�گ_���!Z�l����N<�)p֣��DY*gx�@��r��4?��{�_F��5�e��k�vU����%�X��AD��P�\����R��Jk������Hh{7�̒�=*d&�&a�>�ز��Ɂw1�*��[1Y�!Q�U�K�q-3+�Ⱥh1�(*��B�8���'�ܓc�ߧX���(��,P>"t�SR?�5%���4�i�$�YF�dS���8��)����'��=N���.j�۪�~nHϤ�?���(2"�9��v�H������	m��e@0j ��7�V���[�؅X��b����e�`4��o��+I��v7�U����R����"O��$&A�vu#�Ƽy�MKj��&��!�0x�e*��^�4y]hÚ�c֏J�� d\MsT<"� D��7��u=`r5�Hm0����d�f�:`b�-ӄ��M�-����=;3�2�J_� �k1�¹I�b�����Dwbuk����Q-͒0�r��\���tI�J��eie�W�򤗌��=�
�]G�CK8]\�q�'�"�$Np��o��Vl�v���r*җw�&L?^��٠M_���2��j�B���H�I��ϫ��Ÿ+tl����(#ؐ��e�K{w�Z�M� �曇��wƄ͢ț6�)�#� �;��އ��� ɡ��;�$����v�v?�&Ȥd��N����ufh%7���V�d�Ϧ����r/_�~j���vO�ӊ4Pr��̆#�	{�jҩSYo,x�j�n����N����6`��j�+7�n!��?>�l,�V�N�YF���9�pR�>����8 ���L�����Wr�\���x�_.�1�ř��>�����%{��uh��=�"�[M@����,.ܪ)�$�`���GA��ٶz�?-�3�z�c�<p�;(��O�l��Waȉ�Q�a
񷞐-bC#��g�c���H	��O�Y���"{�����γ��F�Z��|��|�琧�ؙbI(mHT@Ӷ�����o�;͠_���`q�8�nW�,�e#Z�Jw&��K/T�*rA���`zMėg��^��Z�
�u(�������ѓ�Ϛ�9+�R��M��.u	����_��=Nǯ��Pr̥��29��LȮD$�QE�L�N�`�E��{K�lT�t�V��@4�*��E�w)<ԓ�7���yĆvX8_�� �L�,��D�����D�p ��T�S �(��W���ص}����:��S���@(�l��`��u5��0�Z�q�`�p�MBx���x��cx@�Wۏ5W�ȿ��d>9�*�V��P����?���� ]qq�=���"��p�-�Sdơg�k@���7c�*�D��7"׏?O�U����`��ŗ���$��P.R����`�R����#�9�iĞH� W���n�DP/8\��zO��fT:�²�h��r=��Q_�G������J�k��әj�!jfn(�H��l?� S{F�[��Iǲ��ǯZ���˪��R�c6�E��Œ�9�%Ԯ`n]\耡�5��� ,��ˁ~��	�	�
����\2���L}.8�eJ�4�+���U��P.�ہÖ�<(��o������*6��b�~�`��ER�%x5��oXhe��b�K[]n��!�]�1��z��#���]�(�VX�0n�>/�����[f!_��Q?G��t&}��	o�?�#,�3W��}�z��ph���#{���,��aW�P��	��ܘD��0,�s!��ɛ�}2,�8�[z�`�W�FF��q�-|��X5����(quW����C7n-*�����X��\�������p
��L�y8 ���n�A%���P����ˁ��-�$cM��������/�檮���GX�ZC��T�\9�=�M��r��/�W��ԙ��ML��mPv7� �ā�e��%a��5�fV��*�D������'>:��"�'X,a�`.��<A�5PT��h��l���My�3�Q�gzD4���9���	j��=��f� ��uF�;_��9��i~J��(/\&��q�(0a9?b��^�X�g�đ��QV���?���.cE���D<�~����4n<���Ʌ���[,��#+��R5DOȽ�>WɎ�Xx����G˖`5�*�=r[LK�P��L��7��{v�{l榁WZ��@�[�I���-�z_��LF�^��c����`*A���X+Q�'��M�;�LV�~u���NOk��.="A��0��!u�n6�_~b50�YU����$(4���	$e�[����?0fF4C:�D��F���#m�1�n�:�2��4�Ufk�b��H�V��[c�NWE�����O�MS����h��c�ޭJ�x�Ĺ@�kZ��+�"]�:��t#��	�o�q\��)��8���˶3��R�.3M��Ǣ4cI�{C�p���(�2j�!W��P����\�X�<y�5����y_
�(�n�>������qrsM�{O��r �{>�XϬ�A�[���N��F�ڠ��긠�2f���vx�Cz�H��&�+pK�<3�;Rj	?rcV�!�#��ч��ʎ�q?$�!�7y���{��BǬ��g��+�	��姴�n~I6%���hp� S&��ݒvW�?�cJ:-F�l%!'���`EO׬5⁓���e�N��n��~$b$��C���̄����=B[T匥|$��	b��X�MU��!���A��`�صZ�Z����o�lF���k�;Q�*�.�������)=&�*������ W���2ܩ6��\�,��)�.�\��|�u���^"wjx�(��0Z���u>&�D4�"9���np3@me���HJ�{�NT���^@z���f6P���r[4"~t�%��mx)ʰ��m沕z�g�N��5�.��Y��z�����7H�~$a_$����o�6�-���BէM\�����̉x,C�AU� �<��9�k΢e3�g�d_e'(��vG����?%��|e``*�?P��-#R腛���\{�z��T!�9*�4�v�K6Ώ�&���}���ē���⹥����U�E�ָh敾�)R�Rf1�Vaag�\Ip��<�xp/E�t���N��Ķj�����4���3g'�ڦ4��ɀ�<'B���|B��q)Η��Te�h��PY��G&k(��D��<��@����Bd��{���P��F��}�L�ZC-C�3wo��G�H���nCI��g���Ӧ$ ��a�l�U#hR�k�t�]y��b3��g�E�'�-(��=���{;g`:�x�S�9|��&�8;��N�F��a��[{ns����	��S\u�{��yA�w���	I�X�Jwm#=Q��Tze6�U��n���~��p���g^t��3�q`�ƿ���(����;�볼�-l��/���ҝu��E��P�us�J���,�pH|5�����R��Ye&���6|Y�A^w��;Wz��ր�T�!�9�M���3#��:}�!�0�v��AR#�C]�=��K���g�F;X����Z��8u���'�T&�$;��^p�N�]�]ux�%5�4�i��b�T����Ε0�_�E(��vh�if��`�]#� �ߓ�=���'K�0��5s�r���q�Z����U2�� c�� ��<�sW���z�.��B�G����c^�\��4�J@3Ĵ��`HO[���T8D[�4�[٠h�\���2�ws*���l�i��a*1M򱼡�N��������6�\�M��X��y��9ף��1��%A�&��p�E�[^d��:I�SW\��ӷ�llyW0��/ry��\|$��@�?Q-�"�ZP�xk����/3�՝u�ܭO/�3�����b;ۡ���xέ?�˽�T����T�Y��k���|�!P�c�8�}N�^���P�."|�5"�T���ȥ�7��ihS-K}^VJ�B9�a�6����� [8��]�a_g��D�?�S��J�� 4/F[���y��.��r��,�G��p;˟ߖëƶ���UQZ$�ɪ���)uJN�}��:aڝā2h�y�9��J�L�(���*͠�~�C�4���Z.��s$as� #�O�G,Z�O��f@-��f�^�N�x,@�[����n�Ce
���T(`A�:���8\�� !`���B�f^.�xc�p:%Ke��N*0AAp�nҩ�c�j�m��'���3Rp��f��Y|����ź��L�/�.�����ҡ�N�:��$�-���7��I&����7a���mҎ�+œS��0���1E��kK��Ja,��Di���������u!e�������>:)^�+�8Λ��r�����Ưʽ���nQ�R��0��A����ܠ�R���)�Sa;[��S_Y��}�kC�ۃbd�C�5g�����o�~A�gk�ـp��q�M/(3yDF3E=[)BT��������]��U�f���ni&i�iѰ�*6�=���J�E3�H\b�mv�biѝ
���2��v�M`���\�������v�S�c���{�������=�֚#2<rl�J��ocGH�-�n�{����>�ّ�	kx�K3h8�;N��ޘ
~&������2Y�Ꝡ�hک.)���Jږm��;�B+��cg���V�3'�vu�i�I��ӧ��*�(3r\��W\��ā�|NAX�rsF]{�HAq����7��:1O*�P��l��R(u��?P�Q��KF�G���Gy{�G�6H�W��Cs�4�.Yݴ[���V�Թ�u�V$&����%���N&W7?���ZN�&�'���J|�e�H_�l�j�}+7�0A���9&�p�ܒQ�,��h��P3�P����
���1XN����I�@���^�=U5=KZ�ނ�+r�M#����s��VG�v��'Wr���0G�'�˝�R��h���Vm��Q�����cz�����;h��5WwD��+_��6F����g�������d�&$���zX\	:�%7��%�ϗ~����Ұ����YySf!�ُ�S�(� �&�Sf�	ߩ-�� -ՓH���~2��%ah��?s^i��XĜ�bH������hVd�����DX�.��z��UҀ�D��i�S\?�`��p�G���3��Kh�w���S���YM𙳘f�$���o���k��x����#j��:
�j����8V�������&e��'<�2��C�g)Q9�5x�m��g��U��-A��Ͳr�_#i�xyE��_M��Y�%.ہS�M~:�a/�3o�C� ��ou"�U�q`lU�~��K@'�Bn�BA�+�2D�"G3���멧O�{�/�,W��bM���`�4qo��͐lYv�4�B��G�\��9w�K��A��ӏ����:��Q�E�pcA�b���F{|�0��!�Ki��O1����-{��������e��En=�/]�ǈ��z^�I�0CK�z��}2�z՗���}�x�Q�.p�_��eB$U�R9�5��	2�Qt�-K�t����
5dxVb�����n������$	�OpS[s6���=�@j�o��"�)6X�|�~���܇;�;�T�1�h�ք���߷a�}��K�	Qk�օ�q��&6��Swr�����UAnī�R̓��P�.E吜a�Q��D�P�KK%l��8)ĬHZ|��7���ꦑg���ϙq�^!^�*I��`2lB]�؀��§�ϯf3pNZl�.ɠ�����Gȣ�_
ԝ
�(>/�p��u�`7�U��A�+��w-у�]C8�xЈ�O��Ux+]X�-���x�7�z�DE�q���$���H\�嗌�J�qp�H�G�\���` ]H]�c�ț9�i��'� ���������Tf�Lwb�ii�T��ƒ{�(EmC�}�~�Y�B\��Lͼ�+��6k`�h��ĝ!���"�p�M7����v`)K@y�p��y%V���zG��>;S@,M2�S\j�>�,��&��CL����,��C�ʞR�"�ZD���!d�ml7�0|a���p�k�V��n�r7��n&V��!�M2�pq  ?�t@J���R�=�����=,���H�(}���t$���`1��F�,Ň�ĻR�;�^�_&�jVL_H��r2Ey��-R��f�K�J7�S�RA��^*=�eJ�r�/s#�	�(�z�,Ǜ����Zy���TX�d���4אr�GG�)C��62߅�Z7�f����ڃJ'P(��ipl|����N��C�՞JX�[z��t���J�J�ť�.��Wd�x/�Ol ���t..�c-4��L�,��^�����D3
e���f몳$��I��=�;��<�T����j�0I���F�����	�m��W�U/ߖ��7¢i�}�{y� ' TѦ�F�
OG�e��:�5��{j{TE+����G�@_�I�#ً���g?R�� }]i+�8d��w�r��sTF�g��op{Q�y`o]3pH.wJ�M=�׬�zWkE����?#w�R
���K�E�^cc�$g��0�t�@���ˍ*?�Jhn�C��@D���{dX�N�2"��Q+��`}Y�׽�h�z���fA< `KGyw���)Be�+���U�{�~Z�b����f��RU���^�S��K�0�)��*J� �銞�C������M���(#+�a�s:]ua��u(���	�(�b�?	L0A�LII���2
H�'���&�i>�qMd1Q́��@��u�x���.aniU �j��b��<B{ƒ(>��(�?�=ɚ���qN��-:F�_�Ӗ��F�Rg�84̹��fMM��(hf�WG����&ǵ�p���^c��#�a,�����v�@q_î��îpa�M��[w��q��R��A�ur꯻��CD��-��ˠ~�1�:�7E�j,i;v'���Lxi~��;Z�@�����D!�&tOy��zC����gܮ ��C��uՋ�n"����[9Dt!��^i� �O�`{�-�Exa��L[�)��[�:I0�Ũ�����Ao�1�Uip�9�V���[��wj��b��ܕ���g(���g�Ep�v`��,lLAa@-�=I��l-\nzp�J�/bW��á{���-�V�L���U����~�#�8N���}�1m>���4���5���X��p��p3�FSr��%X% _ �I[��R]E���<���SD͈P��$�rJ���x�i�G۔�� ���<���%�U�>�Q1�̸?���9Ȕ�bcJ���n���N�F�q`�^kyG@Na�Q�A>�])yt��]�|�|�j�=A۸o�P^G�Y���u�7��/�J�ۨcZ�?�e䈉_��4�Ѕ~v�I��DQ #٤ѱ�`��Lp��~AȜy�T��C ��t�[h3v�l@��y鳼J��Z�^����-��ĩ/��z��V��;@�N޾7@��n���@dЙ?O)!�E��Zd�V<Ֆ���_Y�p��#�X�J.Sﯣ�s�p���+O�i3~%28�g�� �"*s�i���MU���� b�ʦ������pH��O�YV���ڴ.l�_�g�Y���K��B�jX����su)�
8�T�e�U��h��(Lg�ȅ��GU��;<�;�ī
<@酦��t7<\.�BF�[�D{(�7���+`[��p���˕x�` @p>I�t�'p;��:j�<�WG����U��cwE/w,*g����o�>����vܵq�c.0�Yi���A�h��Y�#��t/�n([��#f����D�24��������h�H.�ӵhI��r0nSe��$߆��C/�Tf��:�2��V��4�f�0n�9��d��w)�x����M���:�?����
L� (i��}a��G-7�Hʡ�?��n.(��v#��ę`����}k<����%6rd����@#��?���d�M$�A	u��򳞀�٪n-�r�^�[R��ʚ[���C���d�Z�'�4�\��،w� {晓��LWca�`8i��s�'C�K��\?c��G�Q��mA��j=�w��_��oKt�}��9B��r�]QI�^��6�x�z~e	@Hc���������A�bkY�8��%�2S������eN*~���r��^��@0�]>��/�{��S�b�����iF՚�ޡSy���G��1eF�,-���b�0�\K�L�r���D|х@�]\G��������w�fƸ�W��>3��|���gȑ��xm0}��t���oLusX�,��4����(i+�(.A����-��A���sZhD;�	�M묙��Oa�i�j��7~}���t̅0^׻�N5;(|��U�S�g�����\C��
A���j:c���Y�:o�Pf�g�2�V�''��ҋ]�/߃�Do(d�l��b\��jT�&�&�7��Բ�֢N�����D��i �Ƈ�_��$ 5��J>��sZ�=�W��N"�J��P¡��{��Scn���o�����3���k_��T\C��y��ES/��ʌ�rob=P0��D��Ӳ��œ�uO�pt��s�6S���vVf�#�"�Ti����I�S�5�5��S�s  Y��\h��א)��hne�X�P��hqa���p����]R�NA`��ʗ��zE��C�*�>�Q*kh�l�X��x=�(B�|��$/���=յ�rw}�F�Aa�����"�w���&��f��|/��/jn�k�Qg�\�B���*7�����՘g0�gX���X�89�m���҂e	9��"3�۹=f�u�ȏڹo�莭5͝��,gи;��/�@o�.F^αh-ݨAv��%��=�����t�V����VT�N����g_�F�]h�������$SPbR�c���b,!�����Q�ۦ�!ܩ�	�?�jґ߼>e�;���5�\�IT���?��â�9��\�̵�.s��#)ڽj'�����)Yz�ǀ*��a�fs���OU#@�_(���+�R^G��	���WB�ܩ��2��
Ӹ���«uՕ��Ź���9���sV��I6=���'�@�d��4!�=.���B�����b�.`�|R� �����ba��jr�'�q�c2K���٥�y�*�u�>Жw��ڶε�p��0��hM�jD�F>��;y�&I�.�2�&x�0��
�H��\�.� *�1I�Z�R�5��!� OW6r�ػv#�.�-r�plO0"��o���m����b��BY��)y�K]���};��ȥzbK�u���:n�6ϝ��o@TT38����_! ��F��iy���E[�9����.Rs��#�8�����%��\����t��rشߩa6�cBȠ�l���K�:Pn\G�<�[� ^ӗ��rx�f�(Lj�؁v���ǒ6�+������@��؋�����T�!%d���x���L�i��)2��q�5Ϥ`<C��*�t@X���M�Z��y`�&�wy�JK��P��	Jީ�

�q���_�fS����k�D?���s6�[���n��O��u&�o�	�����t�'JZ7���"K�*`v��$Vf��>�bQ#񍒰�
Ra�a��ƶ+�zk�lҠ��߅���DX�[���g���Z��DQD����};�fő5�p�uz����&��V�I��W7m\�r�7��iZ�d�ݎ�uC �ҞI�%��%oul��x���q�G�P^�"�<��X�|Am�]ЋCz��@�Z"o@@b��.����.��; a$Lཱི22�pbZa��VV���|�k/�:�A�{+�^�P�ʒ�{�>X`�]O.��!������eJJ�Ѷ�盭��sd@�� ʕ�k�e�� *��)EW�u��46w��!oXձ�n)U(c�e���Wk�3��eaFRi����m3$���;y�����ܲ�q���aC����������b�����:ߞ��є�q��c��H��}��BM3������}�M-p�"W��~2�GV�2��Eǌ�*1}��eb㳽�k�an���r1���M���n{�I��z�V�N���`k�jסwkQ,"z)�����p�^����<n�ˋ�<�H��H��4_n���֋.í6 @��t�bP��/��i�;�i�P���ڥ�Ud.݁��;Z��dۚ�w�R�&��h=��F�Q��E�i� ū�q�p$o/�u������H�vJ,ϟ#j��V(�����[����z�����dt�m��~/G0Zyg�h-��o@�֡���8��m��d2�/xe�M�(e�x3� ��3�-�2o�2�y4`���q �I�v�g�Wbm��u�>K/�8x4�kLR���ޚi��A3߻��l�-���I�Ɍ�Bb����}����j�9XH�o|w��������!�԰�š���q�V��o�aT^�tZ�g�n�Au٘�ge@�(��ԇ^O����c6yo��I��Uv,��\=M������H4e�㔊����=�u���ktx^�1]����N���_vu�iB=6�:��|bN�A���2iN��q��0�WR�Y���%��赕>�߇�3eh�۾TAw�Ayp�:W�l�K.B�੟�� �pdY�Re2��G�+!��1+����K��pպ�Ѷ�̭D7H0s��|`��!6�ڤ��*���%�����-,>���3�z���x�,����V�TCeȱ��3$�&�E�0�>s@u[�����ȯL��ܘ����sy��SwS���F���>d����Df���W��`����;E�Y@Y	��b��]����w�P��w��D�x~���Յv�}@�#��Z1�s�X��i�#Ș��9�Ŀ�Վ~���Z��c���P��y}��=�U���\uK�f��0b� ���i$��!'�[ߙ(�?���;x���\�6�Z�E�tw�8���}<��s�#.��IvS��	��ӹw�����=�o/�\/,׵S���J��IQ�}�oR�a?��Y�S��r�����3����
q߮Z� )�;!r �'%�l�g<p�e������^00���ɟ���C��,��j�xl��6���/g����ѕ��;�$�.A8��S{�"c����;�
��|Y��xi�}��/��y����%ל���%����jЁ?�_�J�g=<�nP�d#� ��i�N[���
�|Q�^���ah��0�ǽ�G�D&�fպ���:��Eͩ~�Q0_�'n��l��?�k��#C��mX�K$=��&pٌ���W��L�)Pm��
w�_�	-B���s��ŝ�2�$��e!_�<�T�ЧU��\��ޚ��B(��:�@E��߫�v��]�Bk<U���w#�c3���W��-�l����,G�@>ߑ��PXQ���i�t����b�0�[a�d�߃�1����*Rs1��[���Zs�D�Օ�@�h�ў�/��SlA�kC�J���i�X������ ��_�LtJI�S�C�ߣ��?��Pշ�%L�{��Љ�My���y�
�	$_Ck5�3_<d������J���`��6_z���>�N���7��{`��/�Wc��[\d�*�#c�Y.��	��zMhX�3S����\��J�1}����9#�XS��7X��#�F�]��bV��N&�h򲧘0�m~�|KU�1bה�V*l��%m�!;�
�P>�X�x=l��J�FYd������ϥH==�zȨ������$V^��M=�*&3� �f��.�{S��Lc�[!.�LN��+q���߽���l��"i[�����/�͛��4/Z�μu��x�B�N1��k	�$X���6�73JW@���!z���x��t�/��e���АΦ�Կҏ$7�0�Jќx�!h��)�AX�Q-��g�q�ZF���.�yc,�����q���Aȡ��I�58����y!�%1c oke-�EtM۟
�B��:]����/���"��@���!{�"��M	5�ߠ�ɪ����E;i�ē>G�u$>R$5�00Ny�o(J+U� ���8�v�y}�9_�����lu��{&��SP5�v��R=YeB"�IX��G��4C=s�K����q-�d���#�'��R�^<��e�iZ��4��d�K	I�RT��\��>#���  3Nx���L���;j��+f�MFx�'O�P�`�;N�ŤR-p3	�8�M�����[�0ɘ�	��৒�@�<J���Z!�8Pﲊf4��˱�/�����.�|k��)��p����P$��YpJ�L3\��f`</��l�}-VM���]t�(�	6�a��!}`�>n�b��h���c�~��/��st�PE���㩼 c���TO�~���j��ش&�ۇ?���g�.\s�!yS��8���6�e�D�&Z�r�?�/�ސ��4��Ds52:�i�B�P��8��z�6�z�Ԉ�J��6"9tq��z�O`5�9x�V,i�"X��9�56��y��*������9�-]�+�L3g�P���zA�5"�DY�H�wԦR �Rb����p������]���4��p��x�	~������S�d(D�2;�*�x𨝂[u�[�|UQ0B�:2�`WsIOU�1�/�}/P��ÿ~��,ul�_���F�֌���䞂{a�g�SN8���=�;��P���[�c����]��۠�'��U"�+�i) ߫Zϡ	�n����<��ͧ/�ٓJj�������K(��D0+��Ir�7��
��ڑi�d	֯+�;X6dx̫,�ΒKx�U��w���
g=��q�ev�ES������ �uCp����)��C%�A����g��5�����vu��c��-��=?�R &ȍի��8�{���#;��=�[��d7����������J�t��2����پ�8 �3Jq_�0m̭�`�|��h`lw��2[���G���_*��-��#�%|��(ѝ\���tʩ\�s��C�̈́��ۃ���Ӷ�-1�2��4�cz��J���W � �D��`��?�A�?������?Pa�I���՗L/"1��#p%���ϩ���Yc�M/��K��<OG�=,?�_ܡ��M��5��:�bCi�����T�����\��Hb��ZN�wr��Ih�]"�>F��4�c2����,�G�\D܃�8�wi���A���\�Ldy���p��O����x�@���ek���(ė54;j�~LmdIQ�����X�5�.f�aqʀ�hn��,Q}����s^*^�mU�W+�6!k�7��e;����~|Q�/oO�]��4%�Q�DT	a�)��[=Oԯy���7a����y�ƒ�X"��/%�e����I��H����x�;��z�0d�cܶjH���'�Y�5��
�H��ag���C1���K
jD�Q�= �?�KݦS-�b�2��<~Ӓ�-�k~e4���:��Tm������\cZ�%j���;6��L�<�_.����Y���K��۬�~�iGc1�$x1�O0�B枩��KDa�l�#��2b;x���0���l�R&4j���hb�?��arU�W�18t�W�}�z�˭�V�3M̌�k�x������*�\,�M���k�X@�'����&¹?:u_�� ��lbJ���(M���0�'|����	�r�(?�R���p�1�*:zVH7ؠt� ����������+���-=t�.BҺ�/���3�K�J&�����R]��N�9�֣܍���M�W� =4ߩZ.�Z��*�{O���=\,��88��/y@�9&m��K@^��>e�4���h�Z�|���@�t�F� ���!f�)�_�]{/;��V+8��0����ţ��O*�8K<������ f����uH�K�Xe|��-����J�]��e�����Λ�(��3R��T���o�Zr��T�q<V�sbգĬK+]L��֊A��G���:|螽�Q��Q �BǮ��m�8{�mO��5M��RF��i��H8z�M87�Տ��ñ��#1D;✛6 �p�6�%�,�N��i�X�f�6�TC[�-�M��#}ă�n,�7]6�Eñ�`��	߮>�#&� ��Nd$̲�F6O�8w�i�J��x�� �q��Ջ��Aqm�>�Rg3��^���lIbg8�u�*��N�2f��x(�O=_��c调���:�h�_<˧���2�ݺ='y���|�C�o.!W�mg�	�+Z_��m��:E��U�Y��W�0Y��*��nӟ�gcz���!��D��=�~�/��>n�r�6��22��@D��N�.t@�d�j��z�=�x3H��y�5�mW��[e!�̖LF�i��T�j�i��Ǿ�\rͅ1�&���FA��F�	:8����-}a��-AI��O�f �z7g�O"���b'�����sKnT��`T���[:�=3�Ns%��+M=0$lp$�D����.;*��!��!��BPZ@a��&�]y����nwNT�I�,s<[�}F�X�8�ta~�l��2���y3L���iSu?�Pz!!��6�g&}�{V�ϳ̖�w�~�4^�2J��(�0O��>��4\��]��Hlp�y�P!�~օ}a"w۱E���u�e��;�"{u���}+��jЯ#S񏹜�Q�����x�\���|`SO�{�|�uk�>H1���c^Z�aZ 0/���,��� �~�)�VN5�+�.�H���Y(`W{�$$��*\��FP1���~e�6���ĝ.��oz���c���b��)G#��w�9:f���Y;#3��c�8�������)�=ŹY5�!�xzlp?>L���"+��Z%߳��1/��'���ś�?�uU�Ѫ���`���d���#$�����ha!��)!e��	�zy+��У���4�N\�ƦN0�8��(����,eL|��+�y1� )Y�zM����o��tǋn� �
b�0��]�����Gϯ��m��Q�6�:m�,�	��>�E-O[��tf����O���wP3�4e��}a0�����yj� x�2��ځ�.�eC������V�lN#:��hw	h��_�e��e�f��;�Չ�ŉ��Mz�w+^j�F;���(���1A�����l:��4�'���Ʌ֢�X�A:�D�o�M�#P/}�y,|�d͂�qc�M��y ڢ��e�ē�u��ÿ��&Q��>Hvt�_�QY��kM��PbE��#���6ڤ	uJ���R��>���rHXʼ`�<��i
�#���\Peth�G���_�d��w�V{���ƌw���I�C����Ԅ����"f�Փ�~C��k�D�r�3<�� �BF*,��zo��!�9�k&E�9W��6^���C�G�U0y+�CiA��� V���W��4�]ӄ��'|;��s.�Ï�J��#)Ui�h�x�-������{�^ͳ�Bׄ�,?-���F�D���k%q�$����
*��Ho����+yX(�D�@�%���K���ΒwV��%Js����+ok�#��5�y��6Μ�
�ьtPV�c��-'��c�s���wdcG���B��~�w���5�c��K#Ԭ�m�:�w����G���j�
?�ێ� 45����䵳;�.�����(��$##_g.��+#Q=K�"o��{h�k=��g���X�&�*+������7����=YEc��C��	�9f��'��{0�����.F�/��B%A��l�u�=I5�.�	�;�Q�^�U��z�!�j��b/�E�C��q�͋Y��f$��"����sSzYQ:v�o�?$�-��L�,���%�]
�^���1�߼�^���`C�zS"����F�7!��6Y�1�ic��5\ŏq�np�[���s+6��F��H�y�H��UUaQ$���<�~�:~q@�Rq�cJM��$��_��*S��О'�Hۦ4��l�|4�t���X��	�	��dy�����<[�:�j�����Z��{4v�D�ؠ���3����Q��)$�'�h�uy�ڶ����9���g���+�*���F�d��p���%��Bg�q�-|0
B��{r�	Eu�f�"I6�G'Ϯc̱�u-Qm�d<�%��K=o�}�Ʒh����DRu�C��G���Y���HE��De̹��p��׋�Q�+��[�E�Z��Z��M�@
��ߣ,Cp]���X/�!��|��UX�mUiglg��N��b��U#,�]Ep��՛�;����"�w�?�`F��S��)#N���r®'���r�\��ڵ�_2�\#܂�թa�U��K�-��F�7�+vs�31�Nx�W`!$=��X��9'W�+5ļ`p�������Jf�*әe���B��y���/�6(�=�N�Kڝn�s<���5�yp�ǏV�H�Qr�A�k���R�*�bi����H=�'5�Lz���P4�+��=����I5�ҧu�Kƚ�YZK��3�
]���G�Y'f�^��<�b�\Pq��~���ԃ+�8�;�7n�??�<U�
�Fh��U��O�T���yzکe���*��#���jM����P�p����,�xv'_S�!C���A���]l����BT��{fѷv�
Q�I��-��XkS�
��F�3���X�� ['�GԾ�bL���}�Ց��w�U*�~��&YLCk�8����{(q0O�� *�oǨ��H�M�����T�9�_�Mj��e�/�p��T�^5��J�o�h��W03QM�0�K�o]���x��#X�l���!	�c��_e������onjc�`;GE�,�<�1ZA��M�f$3~���=X��?h���e�<������KC����>�j��|V�
��J\k�t_:���1is-b䖐`-�O�|6�U��U*��G�r��)�H�.�b�u|1&{(����=7��I�f3���ð�9w,Lb 1�9^�ym+�ݸ��ya";���4L��h·͇:�hsZ��0��NV�G�m<Q��n�ǋ-�%&����bl��'3�Kf�%O�T��c�]*�
8(��:(8��'��ޛ�ΤsխH4ߒ �@�0�O��(@�qR��@�;&`\�	#�:�X��8j�]� �F ``SP��8����2@�f{���R�2�ՠ*ÍF/�}�S������%n�$	���5�1�J����_��]!Ve�u
	�IC�<�	75zfܮ�z�����՗8�'T����1k�E㹯��1�øQ�*�xo��__|�MD�b!�}��ZX۳C"=$�Bi�7D�;N^���,���I�ͺ{�f8�IC�hZ�{s;t6;���0KP1<-y��� �Hw;�IfB+夠-f~&m9��L��8����+�)���e� ���{�~�Ѷ�ĔϪ��W�n���Y��&�oA��S�}��׷d:Ф0y������a'��nf��7X;��j L�C�0��XϷ �]�<'��[10�!,�S�g��7b��4��H�#=����ʧ��"X��V�\
�J��/�\П]�� ���ixj:��}�x-d�|�Ym��9%r>�M �@��*�HA$m6V�IF����Y�l?B�ʠ9۞�hmrd#9�V<"��'0���a6��yNPz8���ݳ3M�5���L8�c_��E��)5��
�ww�mz�5�Lj�_W#�����]\�;���d~���2�c��'�5��͈8�r�Q���a gg��p��?e�hok����$�C֯^���3A2��@�~�|�72�)���Z=k3���Հ�m�͹�Z���>S}=�q $B�� �T�\�QgR]<������k��,��6Y��:�����#���b-��^e����xD����/��ec���?��p������\Q�;Ɩh�˵kƕO*���b�'��'���OW~��D"nF�|Dk&"�b�ٕb�@�Ӕߙ{������`%������aK��\b��*h���Z.��,Dm{��f�������q��S+�a&"J�$��/�ݲ����L���!t���r��ĝ{��N$�uLL+�M�[n�y��&�-��X|q1���7`}2Ŕ�˶w!U��
@�2s����f��f�1ժi8�F�L���=��a�Y��� V��9�e���"3����d��?7����oD7��v �����>�$�"���N��?�r�	>>���BX�D��ߌ�g^� bЭ�`x�l+�Y��~��S�DHCؒ��KՐ�Ū� d`JKJ�[�Y��9b�0�����s'��[z �02�����t7|Xk1�&�Ue�@��^UAo������R*�;e�c�����H�"��J=�7XEE@X���+�#��8�U��V��f�g�᝵pq(�.�4�1qd|D$[g���l�u;�ZP������
STM� J>�Z���w��Vc��x�RK??��#9��x�������{d�\��>��k�"�_���d�&��$M�$D�h���/�s�h|�PLX �VQk�.�3��v�.��%l��X��@��]� }�b�H�Vϲ'E1��:(TX#��=x��a����U��PM�oz�s�����+)�_k#��G*fz��"(G����?�K��+9����("�^#�x�(��庰yYe����4��Ue��
[�蝞%y "+�5������e�G�}��k:3�Q_�jw*�*`OX����j�z�5gy`x�HRۈ�����6f$���Ѯ�'!��%dT��!$!V�W:��GU�ʧR�j�:vZ��>�t���F?'J�w�V M*-��K�Ԯ�*��� �dQ���d��o+�d�dVʠ��q�dΜ$�&lTH�큦�t�����[� u�YK���ؓ��3!-����kfn6��!�x��o��%e2�}$ Zb�I�M��|@��g����yjL��|z���d�Rݳzx���������E�A��N����x�ܕa�(�[���H���q"�$�{3/Y�>0��i��ug�u��5�;�W{B7 ���B�.���z<u�î#�o{3k)=ǧ���ӯ�S���V��2z��a/�`�3
��A:��[)�u]����fzcTJ�O���	�[F�Fz8A4ňsA�H��� �2���EbC.�����n�P��Ob�.��X�'�褺��tw�ݎ	�!枉~�^�+F�kwƋ��}0P~��5B1 ��E<��{��(D@�[�;,�9|�VF��P�XcC��C��i�C��r}�ڦZN�^pX���+%�{M�^�<n	Nj1�������������f���r!�ll�X�i�E��dE]����b!��o��0����x��[�_͐�2���).�Q�O��"\��6�Xn&�H�GU_��E�B+��x;��3Ex�o{��wq���y�kd���X��޵!�WN ��4�xb?��x}<@��q�A��]K��5�Wщ��yJpA\�U�ix�蚚��qg,du�<5��Xp�|���g��H����)lO�)�e��l��A�h�iqe��l:���9[I�W���ZH�+�Rl��;H�O$�.Z���W�"8K��w�l��?ja��)�Do?�L"�}Ub���Xtq��� �����\LW�Q��|`�s��.��uQ\�`j�_J�_��TNO��/�3�=�*i8�h͆����m��$_���!"�r��pJ��%V>��^� n������V�A,0�`�V��O�˳��b��iF�>l`˟j���^�Q���JN"A�%Wy�d��F�V���Wʏ��\��3��%�Ւ�	Q1�b׿a}aW�D��Q\H�F>�LqnF0K�ђg1^雓E��_z~'��Km>)���࿬9,/#G)�E���ro��^c0�ӯb�(��.i]�h3wSs�)���''E�9�>mb��c(}�6C@2�@q����Z�!��=Hե��s1m�M�Z�����OnV��)|���?K@�(=��Y7�4����˚�.�,; ����ٽ�vĪQ�M�V��(��?���U�ei.�>���BS��V<�DF-����|�
v�zò���>T`�'qLN�=њ]��PٵƑ��H��NB�fnpʶ�v��.��O]�{��qQ�?��N�: ��J�@&�0G�L�<����<.vq|V�TeYƵG�Q)�H����l	J��g����Tu�KB�i��ߪ��	U",�����#y�Fr/q�{�33z?�Ś���D���Iɴ�2�f�i@���ќ�*��y�j#13-�G���G�}�]����.�ޮ�3�*�W6���h����
���j+�r`b~fZ87i5�:7L��� %!emMq�E:9Y��uM�Q���ŇV�Љ_"�m�52��<���@�?��xa.����i�W��J-���)��4��>�(k�0�Bl���z!�6�}���3�o߬���Րz��O\�������;M�Y�����OG֯�/��g�|]q�T�x���k�u�Mt���H��rw%�^-���i�� Ɉ���9����Y�_��ę?%�*o
a8DPb��Nl��`e��lf�kc���=���#;1�ͣ��ڹG2��ٟ����=~��Bg��������dl&�� �ab����<Q�ʤRmj
�=���L-�u�3/ϲ��vW:Y�z�������a��?�Y�� ���p^�33Z�����H߂� ���&�-t _z.�4��(�!����ދ��tEɌ��d��=���G��y���,'��	���x�����@��ȏ�I�}y #@���� ,5^;[���r0OX�Ky||ěC^�&�dS��>�cv>8�"4��X(��Y���aF�Fv�mE��´2VZ��l�kM��s�uǅ#��7�����H̪&�z�t�2yP`ል2YM����9�=x�gb%���y1��6�@WX��# �sE3!:i�\���5^ġU������KT�e7�P��۩�R�"ڴ�&(M���8q�W!��b�E4�?������[ɻr ҈#c$9�<�Hl4�yi�r��a����U*��.=�M-�'W{�����;�^5"�2�OKǊ5ɱTfѦ��r6��!��S����2q�#�I(����w�e|,�b42:��k~�O�veM��Ɍ����[B��=
�-�Q�"'�N����2���2!z���)��;��S�������2qc��@�W��vPN~�R��L��0��,Zsf��3�V���lh<�;6N�bQ����YO��XZ�l�b�{��ɆVl㌈��$�Ф��i"���-�>�[.Ŵ�H7hNv�b�B�t��Q�i>x��Ѥ��C ���e%��|b:OA�đ��&R!�r�A}z�0\�*��-vC�.JB��n{�[��ŏ����jq��!�����[P�HR��H0�">��ɾ��E�^�z�f���$l�˳V�����C�K��kZ�qލY�������u)��1�z�w4%��X_VN��{+�K?�Y�^��H}1�JA���<�u1O�	6CFT��p��{.()� x����-R0�Rݰ��5*N��`9p��'�/�L�.d>�6���d����g2E3QZ<R�;X�?���)�`59|O�����s��Τ&
٣:��X����� �|�m���l�I��+�˾��#�ed}�@s�o܅lTi�!w%�_��I��Id�=.N"��z����R�LȖ���� F�]8�� vӤ{ڱ��%@��j�F�s*�PZ<���_}�=���rT䚗��C�0�D��u"�����1��,����L]蚋-"O�@����E^W�uj��������z<�ü�I?�{c$��%]
:8�	�ٽ3��^�獥*�1��{�'F�3?Ģ�]�=R]��$���^����z�r]Y`�uEF��� �����=ϕ�������/�?�ۆ��5�1��g���]�\u{r���Rw��_5�֨��R\��Oa{���d�j馟z����Z�ײ���=�(��O�[��c$�e�&=*�[��U���|as��x���u�Iiz�y�+�a���hm���;��>�����1�}���L�D��`ar&\V}�P�p�Lo�_��aDk'/X�s~����<@�-E6El��Z�k�̜�� ���*ɀ	:��=X#He�J�!	��p���q����QY-���.*r<y�y�n��A�!� {ƍ���n���m��;Og�b
��k�	Z9,���W���N�%��V�vU7�u�H����@�t�x�XҸ)5V�kQ&:�X'��������������4�{d�cjdT�T�qK{<?K@7��=
ě�	�\��Fݔ��������<E�[4g�����K��b�ԎT"�u&zC�����I5�������T�L�(���Ā�Ғ���D�(Ex5���ei�
PEHk�`�°!in���t9�9b�~����T�ܿ�T7��c��~��̓/?�,�%q������<�X���k��\Q;���a�*~ɫk���#��h��lZ�u��/e�&O��Zq�}��H�n_��C[��(ߵ_é�ڻ+ȞO�JzIq�s��x[�U *Y���Q�t5 ��<��n�%�5g�wf���ڛ`<z�]v��Y�X�]k(`�*�Δ��J�{$Ч����?%"�����I�u�=֌�L5&3�� �k���`j)-��Hu��
�E[��y~fh�'�����m&�ՠq�F��ǻ���������f�]�}�.�v�4��"a��!S�����VJ�V���T8@DWP�|Vӓ:D���ȇ���đ1?|�� �.�y�'�qӫI1GS�9��(�^)R#vN��r��n醾��G!?�
����%��\���� Q�%���)���XFǧ�F/26QNt�����%�8�w���M4����<�lȠ�ƍ�!TO,9`TN�JMm����ÿχ��{?��V&5�VC�| k�2_���)pxK�J���mLS���e�����y�6��v���ǩ����UĀ��n�7 �����H���hʨϋ\pgI}���jUQ%f*��J���F�	�s��}���vO�5]�iZ�2Ť�fkCd.
�gMVі�����CO;���zS������p������M2��G��	{7%�;0;Z���vг��m�	]G���,��Q1<�c�B���p���f'�!v��q,ڧKړ&OW�a ���6�Z��A��2�F|�;;NGb�/y�k�1�94U�d������s��?7V�'Џ�K�p@W���x���aŦ3KsC���{���oc`aW̖)�^���ʇmi<��>�-��\WI�y���A}��5H�����0n-og ��?=���®a>I���S��J��������2���x[s�������8~n���6�^��=�濾;dIA��y㮋���@%D� ^��_�]
��!������X��B������K@/JTF"	�N�ؑ�h��Пs�$���b�Ly��@���@�_J�� yD�n{�yA���DZ��)�SQ��{�',��oH,�^��&z�1���LW��Oӝ� ����1��W��YD�I�~�)��6��L��>T(��q/`$9_��Yϵ�j���;}��}������s���u�Uu����2e����"���@R���X�d�^pc����6�wU�񚔖EO�荥;������t4ʘawe�eڀ��!����<(m����|8$��:��K��b�=Һ8�x4�"ꉭ�F4�c0Mʽ���v����+QHk$��&���7+���gg�<�Ӈo!'\�4���ޟ<��E��ԶЏ�_�����5�*�B�� ��C�L������tN=t5-N߽{h0
=!dQ����L�g���զ-�A~�Y�ǯֲ\��;�`���ձ���^<�n�ؑ�d��
1��w�WE�v
���]X��tMO�����w�����r#�26z4��x�WR;Qu�_n�v8X��8�ӁZ���'?<��6#۸��iA��ׄ�u��>��&F@�~�}��3?<h=�u���ǼQ��n��w���gr���6����l���J�������vc�J�9�덪k|t���Hi�X�-���1�cэlP��|�y��5�JY��u��o~��I�Uږ����Z�W9�c�ܾ�^N�g��[$0�<g��� .��R�X������g6M��˶���x6�h�Q�w�8 �p�`�Z�)|ƒ�0�`������ү++�7��Xc;�����}��I!!�U5�E/��f����1%D�n�d�Jw��8��F��qJ�����|�.��� �km��$�/�UԠ>�9��>_����:����PE�P�#�&�r/�u]��K��p�D��R��i����c���l�.��![f���ssO��#�0�3�A�`V��-as,�w�]�\�p�3�2K��QSRn_�� ��;�%ZJ�X�07�&K%c���r������@���a��ۖop��~���l����Ծ ����+��Z��-�*7����_�":�ਖ਼JY��VI�ƘJ��ԃ�,&M�̝w��o:�9%UQٖ@-"��0t\�\��a��}j��]��W`b�;�z��ǒ���jRT̟���͔�2·-5�����'��Շ��G�f0����`�y'�Z�!���GS�,$)R���Z��ܠz��y��H�	�Fi��6�=ѷT1O������wD/`� inp�$��PkkV�4sW��_z�S��L�i����H�7j!1�(�f3 ���On�F�Gkw�^�y	����Q)a���#��E��9������oto�^`�3^�ց[;� �0�}I"��*��)`}���3��y���s!� �4�h��]����&��\Og��r����@%q2��6Cδ0*�]j�Sў/7ᴳ[i��X�R�`N ��m�
9N^���nnn�߱�t�(�	,��*_�@�Y4xvR%x��3����R�^��(g�+V����OTa���W8��Sx�7��[�ۓ��l|��S��7�f����E���o�^5"œ��8�?�O���%��\N�Χ7���b�6� �MB�l��H>����nKݾ�>���G{�򱎜��[��vpj�����F��}]y�h+ٳw�X�ܐ�Ю�0����"ho�����Y���"!d1VOWa�Xa��+a����S�G���-.^xJ���$Gf�TcI���|�d%Zp�n�`�����;�+���,s���e���5�0�`q��Y%f٦m;��#&�h�$`��5�����Ԯ��ߤ^��U0H���fJM�R�d�ch�����B�WA[�xE��Od�~�]+-W�q)��0!V
�(hw�Z�B��إM���#�$B���b"��&����+���YEc�դ[ғ�l`�Ej&m-�;�Tb_l[��������θG���"5��s�#C@��B��(m%����b:^�^|��s;E�r�a�9��k�J�?��uX�mr�5����)���"�p�nAZ��{����9�mu_�١��G��w�Q�,:IOvo9'���ʹF�ɻ�� +��؃�U!lY}H�l/]r �4�2�� ����N���MF��lDuY.�r��KWr67*v��T�6�v=(r:9�jP��`��Ŀkm�m:Z�"FA�{���Y�����+�j���+�Ш�~�����T���#�����!P�J���B/]p��@!�i�%�fev�7�>Rߠ��Yxi"j�%ΐ�-�$�u�x�ެhGt�nא���v�Rd�҄nmcܘ2��Oz\0��0�#�b�J״p��O@�5f�����>˨���_s�]w|o�ti� %�^�M���~/���Gx��a�&��0�a�jz�����r_aK���Ygƶi��ȵ��r������|.�ၥg��;Ɗ���f�x�7���Č�1u`��j�K��fE�8������R~(�v��#n���y���ZC���~�2 ����zG�������r�h|�q_������!l�Y�z)�[��2�*���O}�	���ڢ��0ھ� 3�c�j�D���Ȑ�B����Rΰ�W�����,I���Uw�7��������1)�JD�bn	v�u����RZR��Oų���+��9����V@+Je9v�vˬG#�����+ϧ��QX��j��S�%8\ݎ�)΋��W��m�W��Jȑ�1��x����������$P�C�j�R��J`�2de����l��]�[�.[:Mɰ&uyX��GA��AMw+�<�����aYYs�S�F*2�cj�e���yϔe0@����K��0�4�+mo�x��S�v�ăA�\q�k�ycr��d��(O����C�c4�T��	���1^��BD���i!I���%����˕A��$k3wI%i=a��$tE�Ǭ�\��F/!j�[�FI�F`�0�q�#3ο�(����e����uM�!�?Y�8(����`�a|�2ө!�C������#�(ЙFH��/W�����v>m����;m��ѯ���Ey�iPU�O�Σ;�2���kǈ~�ر��Zn9�S�	ڈ��@|.#� =��E�c'(�ҍ�J}2mxɶ�����Cc��	:�=U�Yɖtb��O�&��BU��n�hġw�G��)�T9S0-_�3=:�`�rX�k�Z��/%}K����y�o�s�*O�0/�}���DZ�("���Fx�i�|��u(�˓31� *b�9���)�b�NxU�C��}C���A��D���Z�0��+�T0���B%`���t����.�Ы�R��σ������l!�@��V��翺O�\G��!Ġ��B|;���Z�۴/�T�hjG0\D�y!�3B4J�3-�(a����n�ӽB��gy��A�!$!�!�v�S#P�#Z�Q��0ΧԻ��(�NM�{.tR�b����V�ȭʀ*�P��r�M���S���B�Y��@�1�C�x�ԎR�(t��YS���������~@P���,uznQ�0�#���2BEX�D2�qc�(�� =53.S��`3�V���>h2��~_3�v��p�y��s���4�o)��&�~��2Q�}�j��y�J���3V�EPK�H~@<� �%���+�1�fZT$x�_p{>�`4��4�"Y\%�'�VC�K�0�*��8}J��Sŗ�h����.\n�2=�O0���)2B0�����$�b Xx�j7����t75!�]M���&���ޛ	o��v=TJ��Xc��$�A��ޏh9f�r�b����u�ѭxq�ʟ����<��r�yYɫO�5�����%�t�
$��1��Ǎ箎d�zL�o53�1e  �i��1UI�� '#��܊��=�`���E�!��]�ɱ'-���~�'q���ϖ�����(���̙8*��(��p���p�+]H4�"���y��,D�<?��͑>e�e����vG��8R;��I��aWd�_X�EY#ٹ�z��A�t��d6����N�đS��KH�צz�3qnyüq�(���7��jɰ�ye��,��a�658�c�C�`޳r�Z<hŏI�猗���C��q��������F��F�9�b�]2Fj�:l	���P}#5��6v���Ҿk���T�q,�3��.�	W�XǸ��j�sr��� �e��փ2R8�{pV� &?PȒ��~#ҍ��T����,����+q;����U�O���*`��g�8�q�`��)���1����z�)M�t�yKH��I%U�������;M�<K�=��)	����cky�A%�Cȳ��>;�����S��d[�"N?��w�;�tOP/Z�[��#��� Xp,�����wݱ̶㺚a�w���t~1�>����"KՍ
���d�n��J���mU �����.��G����'���t�GV��{�QG���Uc|�;���ia���d:<0��3B���}a�ֳ�F�HB���s=��N>p-�;��H,�Pg�8ص3��va���ɻ:��`hecX� �2���J&W�M��o� �3��p�!N�	qeգ0���$q���>?4um�&4��t�T��J�@"�<:�~<�e����"xe-�X����VCp� �a�1���7}`�x��2�u��dc�c���hn��9�@�Z�t1z:b�/������<2�R�h��\O�+7����3Y�2�t�y|���.��ڈG����"�N���H�V�Xb$m�-t����~ΐ�rX��,-��Y��y]����b�̌l�\�Ȱq�CHJK΄TQ�����xaj�8d�z@��іO\��
S>rU��KO&����P�7�`Nؿ���L6<1���N�]*e%h~D���a9�B1��oP�4�NSÔƬJ��.���n3�qб@3+����Q�]AX#���/�����ګ:aD�u�irY?D��[�|ŧt�ا�T��!~HL�!h�_ uօyBg%����V�S�:�	\������k�Y;�oif��'Ž�+��SU�U~ ԍy�, �2���0*x�� 6L�<mI�W�I�}�"��+���q�A��%��x9��[>u�˒Y�[�=^:j�K�5��A}�+�h�X^��v�)/�E�Ptu��S��d�t�D�}��c+À���Ѭ���.$�Rh��LM&^+>.<��GP;f�e�_la�)��Q/���&�>��2,�b��["���D�� F��z�hhf���8�G��� m�R0,�p���)��|�+8��7)3������ъ�;8�l�\���1N ��w�w7�p+/QvwP����j��ܣpm�D"����ڏ�N\�5]�K�;8?J亲�O�]#4 ~z�z$��3 /�g ��!1�y�nm�X&[�*F��u�;���
/����X5Ʊ�KSo�h�o9�'2x����6���J�%-�U��>�R�pY�O�~et�}��i2t��p�ae3]iA��hr3��_��";d�U���)�[wm��7�|��#��gH%Y��=4M��G���j.��t�4���L���{��Ur��6��Z3��p�/�[>U@g_�N��O��{7Q�w���A/�f������'�-�5�C�_Kb�����{1Rs��R�;���0F��@OBW3(�#�E�|
X��J�-fx��MՍL()C��z�u�ai�q=ZʏW�X�!��y� Q3<�▷�k1�JL��F��������]y���s�a��	bK7s4EHM;E�\j̀fEK�B�V��7c�	�כ�(�'�WU�F�����yD�����9��!�e}k;x�g����
w�r�b��2�e:������f���j�4q������"��K�w�Kҝa�X��Gł3Ҿ	B�Hh��H��1�\�Ԓ�G-�� ��e�۵�� f�s����&v��AQ'b�s��uM	@t؝�w��~ظ�v5�]��k�>%jF4�kB{}�]�$��'�kx�\� �i6p �][�q!�顦�õ��������a�:^�j���t�9G�J�2m��0d�W>$��b�c�s���������#@w���R�N���mߝg�e5x��燸������
�}�$���P���h㚌V�-&���}��hW9�hk��U�p�i�c�P�e�P����G�(k�ƥ�&��[(3��d���ܙEa��N3���en�µ�)0��_5ϩ�"���-2:��DN�2����w��}�+S(	މ�5.=j��_D�1���`��͈ߖ����X"�2;$��F�]��V�ϗ��IeG˫<���u���<�`�q�t�Z�5Ij����r�\��-�1'o|jW� 8��o��ѣGz�B��������7�)<����f
L:�[���u^��6��s򃞃5��|����:/D20�I3���I�qP��J{��J��}df���O�$f��?ir�����]������Z~G�!��|�� |t��AU��"�o&���4��Dbs?�b����[��=�3�����k<�@�bp����nw�GzT�܅u���\�5ላ�赎�b�W&4]|w{�V����o,Az�rw�xd���{�G�\ k`-��hM�ئ�&�5/pyD�pd�� �1u��V�?��b(�{���������;S�6��s��y/0�k���py΂["7c=Op��B����!�,\�I^5QM��f�I�j��w�ӄ�I���b������("�NmJ�x�tܕ�L�Ly,���ɑr.�{h(�l�-�S�-^��=Wװ	�.�w���G����j� ��{onwǾZC2�rF�,�T4n]��SE�ׄ���Ws�}��J�L�h�p�;l��a!`/�J��6@��y�A��J<4�LT�I�����~�9����V[�Lp|\s=�m&��[ԏ�z�����Ӕe�i?L���:ƅ��4\F�	ٚ
��Z��t�z��I g�*2�^�?3�Ye����[^h�w��9-o���+��Y6l�9�b� �����z�h�s���v��� p����5�6�h���hᇍCţ�/&����2j��]�o��La�ߡ����(�ݬH����t�u���̱b���Ξ�&�GIi�}���@Q��pu#���B�l��)��"��'�D�D��k���,�i��5���^���4��-�p'	P��%+�,Nź$����C�4�f6Q�&�g~���"�p�0��v@Ѕ�??ԫ��<�.�{���L����]Ð�%{���.&d��U���w�Z&�t��ľ�� &�5c1�*R^c��6�>ޅK`��v���8��Y��a�ρ�&�!<|͘S��%�3�ˡ�QLW��b�L��� �2���8�ڊ�Yҩ��}����܅���e����b[�u�����R}����Z��Yi�Q@�R^2I^�2��)�+���.|�2/�3��)�Q�[�wGN%rg��|S�:�+Ź7H�?gN� 
��P"���	W��ӑU�%uha���i�&׾�LϪ>��z iKk�R�
�[�z�x�pz-ۀ�B�&H~�b���C$ݖ�$B�Zk��\Yp��b�v�Y��IM]R�]��Q��1H8�����g���_���p�]�������<W��p����#���^�x�j�U�n��p�"�^�4PN�D̢����y-/�Fm=��?��HlUM�'Q��-­��I�~
h5��Y�c��({S@=54a�����˝��k���*�cf��)42Bh�����K�y�?���O�+��OW�h��_�؋b*�'\�~�V����؍��)���o�+��p�.�Ξ�
s����/8s��*� �_��n#=��3w�J�b(��(���1��Me�R|�"���m���ǿ};��u��Z[�>�D0�1����H��e���wz�,zu[�)�[J���͢�O�{2�{�@�PW%�sm���ge���B��D�2�O,��R�;�/¸��*�1]�����Иw�p��5�:@��@�R;K��XG1z���ae�-(Dm,�r��E{�/��XUŉP�Y>��ڊ�@ց���p��ZtQ�g����V��|3�H���X�ɛ�ܯ���W�g�=E��	�uZ�-w$�b�J/E �~Fmָ�G����R��-G�`�2d�ӆ!�d�l�1�]�#r�1��W�w
��&�i������$!ߥ�k鮙�N�i�r�]m��[L��W�ф������<1�n����){>�Ѐ(��ʖ���\�F{�u�����^a��а�g����]KjB�atY��-f��ҳ��T�\xΚ�2{	�=�	`|�������9(��x;._Y?J��kYG��� �U�r�<o�X���:�'�Ӫ��B�zf�.C 9�:z�0�.���JsFm�����xMUZ�|���,Q�@)F����6�{���2m��Ԇ��h|�2����1Zp�SF!�xJɼ�|�}�j�w�5�q����)Z�2}�࢒EN��-��'�i��I!v�p<K�l��	��.(�?��2�A���d��ӚEW1��sќ�01(y��и�DP=���ϗ?�V�w�}^���%����nY�O,���t���8��WL�?}��u�aM�E�8���i���wa��A��g~ť����T�
��Y��1gB��Zx�"�ï�D�p9�6�2E��l�獑PI�e�?��wP�4�r���������i
� ,xd�%�/~����HC���I�u��p�����s��Q���ߠg�k��%/����MaְF�Dn�!ufY�V<���7�� �����8�{z�,|GpÄ{��Ѱ����8�
�9��1F�=��"٩�c���RĤ��.X��Λ��y��sy������Z�q�o|g�q	!��6R����ߔg]B
��.VM^ޓG�}:7v5�D-�Т����l���:�%%ㅐ@���BR��-6��������w�u��z��	贯<��QO�3�NU����Կ�S1� ؈1�bݐ-�]#̲W!��9z�\�˩�u_�GU�CG\���y��q�y@@�Q��W�Q]�t���xH��k�51y�AT��a�G*�J��Vc�#'���*���E�͖̣��8���IĦ�L<�t��5�� �>�Kb%�k���w1����)�f�3�1B�vp�+[v���z��Rx�[�0J�xh�i�Y��bi�V��69�y����C��fV�^e�w���5>B�57/nM�~]����,��4l� �J�s/,�Ǻ=���_0��S^���D�h�:8�v)�Vt�����<�U��i��\��!�v���������7X5�\���s]Ds&zT�R��`����u9$-+�y��Zl��`����b�Ƅ�/2c���C#����m&Q}Z����0Ii�O�[��M�W!VMR�������v�w�r��r�a� gD��}�qì������A7�Rp�������E����L}���>����m	��/����6�$��N�-NO㳓�\q��nj<X�������,�4�a����k�W<+�
v�~e�J��`�b*��Cr��(.<�5q����Ƴ�^״�w�³5��,�(R{���2�^,���9�V=WMt����%|Z+�j�>,6ڨ�*�\���j�b��FR�DX^��|�f^�C����D��$F�|ГҡX�O�x���^���T:j���dƧ��BNl^�%̏��rg�I���gM�xt���p�u:7�?I�U:����2d�e��
� m��(��R��
ۤ��$�]v�v���i���+�3Qw�Ƌ�`+�{�L�A��YߥE}����R E �H{&�0�/�$?vH�#�U:=9CUK�_�Ǎn��7ȟ_�-}��k�<�Pdg���L�a9�Q��mt�f�eI~e��]_�$���ymը��]��_�P-z���WkLTi|�:̓��v��w��kX9�� �hA1������Z[���v�<B���4<�񢥰��!9`�m�~6�j� �̺�;�80��&X��89;�\�>�Q��B�QW�$�W(����$hR|/��ފ-n#�=DD�|.c�dSϲ9�嬺�^��0�.�(��R�Z���Q�-h���E��p�J���l)��bsŵs�1�].ʷ��+k��'bKȓ���ӳS��!6���a!7� y��(<+R�[�%o�0�g��U���0��i|�!��W���_��*v������jݓ�U
#o��� Ҝȯ��~�[δ��$��.iᙰ�3Vex�RKy!��>UJ�Dx��U���`�X{�y�rL-��^�։LʻW�tP	X�@��3/��=��B`��������������ZOC���пX`�8=��E�'{M�A��Ʊ������i������k0�x�I��oV*嬣��U4�n��1�L�L8S�cd��A1����X�q3�I��@Q$�V�[MZ��Ԕ�J�?B�gu[�?oi&�y^���ɋO�d���q�,Z �ZYH�J*��9�����z�!���K����n��-�<�C�o4�}ޞM$�֒0~���V:�4�:�(겜�͢��_R�h�?�6�ؐq�&�����
����ґ�)t͍��"x��!�`���Ll�`�g�G�������?u���[ �Y���Bj��(
%���j��ɶT���#�?-������H�E�"c|]M�B�+h󚵹	x�[F@]�VR(|�>�qS7Y}��#�����^��x���Ĉ��Ǚ�(	����-��_�hm��.� �z�w�J�fT���f�W�8�&&�� ��Q7l&��!���WM��Ǒ�/�`��F�$bT�jB�c'zݎ�� 
����⌶^�oY�g~{�H������=��!���F'Is�CS+X����lTZ�NW����q���ϊ��ߠ��挾Z�5���F�>���Ǆ�圠W��2�H��P�'�@�6͘e˒��k���:�D���S��j@"�?_)gHh�է�B�}}���7�x.���Zj�f�[P�P"�#�i~�9	FzL�-�3.@�i�	�>O=ռw�H�2�jUzji~����~�y�_Mc��|��ﳝQr\t2q�{@����Վ��tw��'�s�R����뭋�l�+�u�����AP�?��|�����mJd�m�oHN�-�oL4
L���C5�.�:j,QBq]͖�M���B��̖R�ه��<o�͆���.����IOK;���y�x���2��+Eː�`�3��&HR�ؤRP6�ʥ4���(Bd9�i��uW-��)�P+��{i3G���:҂ZK.[A��`䈌�"-V�G�i#F���X3>��h�]u���4�ɑ
Yq�H&:l(�Y9��?�_cj��|��V$&G7�P�`n�%P'�H>g5�@����I�A#\��Oq��	���$�e��)\Z��<��Pa�Wb��n,���d�2N�t��+Q�:D*�Y�s��pQ��8J��Uf���|q��V> ��ŲܻH�T]�/�Cl���"#��z��Bb�3eM�
>^}�$���_ѕ���N��x�os�fIP���J���*J�{��9��I
�gT�������Su6�J]I�BVx�""Y�A�o
�xx�w���Le@ą������r��]�m�:[���b~&[@B��Ϸ�&����id+ߕҔ�#o'���B@@�L�+ې�ec�QlWt���!�}���`\FIrU/�V�X`!��Z�p��-K���*��[ �6��. 2܎�I�(��ĥgU����*���4&�R�&rz�i[�m�,Ovܳ������j�QS=�)�2dwء��Vy+6,z�iFלl3V
t�J��4Q�7�� h�VI���0�q�n��/'lm��*.aҘ6ր%R�j��H�!I ,��4�Z���t3�A��2�#���E���m�#��cW��ӹ��#9?�)�>-S�\��;&��[~3UmO�Czv�#�2�?�Y�)y��Faq�/��v�Est�.�k]���)�GwT\O�ꈃ^7mxq(��q@6��<�0��e���$���Rf���/~����R,T��y��@�!�@���t���
LU��\�N��N\�]�<�l� c�����0�\�ugo�ɂ��\ƌHlbd�C�ޡy	�8�!�9� �:������*���P��U)ׯ��ވҴS����!��%
+�l�*��6�}r��I��Y��F$�� , ��l�m�S�1c���ȹJ�g���E�t�)g��zW�Y���QB~o��lZ�y��G��ӟ
Fm����vx=R�W��ȍ��eJ,᭣�$A��Hlx�C��}��Z���#;;�ī'�EO�U�U�t������'��>I�R�i�2|Cd�&�H%�
�׆=7ݶ�e���w*~�<��u���;�_e0�/#�3GIp��1�o�x�W�����A�}��G���Y��~^֎ї���bW����z{*";�	(��⡇���Y`;m]5��HJ�뻿�����\�m�@����_�Y��Nk��{m���;/;������ZcjM�䁹`��)KVe%p������P�.���c�&����?���:��D�Zk�lV[�mźQm�w5�G��/�~ߑd��"�=�L���IV���L�W�>�	vj����-�nn���J��{�����I��U������h�1���B<��%��PTqs����C�c/�"���#�kٖ�S��DY��Cv(L�-�~��,�Z"��G+�V{>�	"6�u]��=	��ġ�xYc�ip�����l+c�ǋ�Q��4*�MPU�0�T	M�3�i�J3,�%�Rd$�8��\�[�o~=�����mx�[�'�rG0���<LĂ�荕mRh��1�l��(Yf��]������s�q���.�`�K���I�F��]����;�Pv/f���<��������� ��d|)]غ?�!_F�AEA^/CF �}��+�3`3ǦL�� S��%A����3�q\�==[*3^5 �v�"�pWf}#��a��"Aq੝Yav�t�̵t�K ء�(��+�=�D���������������DF�O�ܪjc��zs
!wA��kl�U�f�8,I�9�h��ЇeNz7�M��n�!�qz��d��_��f��Z���Ͱx�RX�?��6H�9�m9��IV��/�&���M�J���~��>�ݽ�>0$�M��ŧ=�"���V~�&��˨p�t	xue��Ɩf�<<�r�xES�1v�����j'�X7�����}���ԩ���H�rB��~ކ�o,ܣ��2�M����z(��\+�+{.���S�H���b������!��	���G�}�ӣ��g�k ��cŉX  7�T�)���,�kF�\���]�xZ}^��W�^����iFԭO;�g?�����h��	{'�rL`j,�����b^�R� �~�t�"��?��O�~�2+��,JK�Ϣ�>}�u���߮� � 1Ũֱ�y��G�b�ƍW��:�� fd�;�h�M�K�)8�]��
:�f�PY�c�������֔�!6+�>&�!�Am($=�Gf��{�\�z�4�9�\����̎S�F�׍���s"��3���T��>S.�a���OƋ�i��#`�f�7ga%	TEZ���S:ă(�&d�+}�n_�뫘�������ND�i]{Qxc���%��"v�5��*뛦�.l���bx����s����˚7-|�Q��a���iB�D���(=m90p�M�
�,��3�bʤ���ۛ�)�h7�
 qص�>�A�`�g%�0���M���<���aT�d���r�iMP~pk_2f`3>٩�@G#�
M��(��1���)�8B2���i���0jx�v��XζA��ۮ(��F�иa��ۧ77�QM��b7�Nĉ����j{�x�܄2>xq�A,����Ϛ�S��-TZz(�'QG7~Zᬃ��N�Y�.���+W]
&_f)a���-���`)�B�����l"��-�>���w��:Ϣ��߯�>��_k6��譄w9�rB�wW�L�|2�8P`�B�n�vh�v��܄-]A������S�[�lt���d�+�exr�ъOh	���/�'���3���\U���Q��
J��>P��Y�Q�s�����cQn����#c�RQҹ�Ϲ�o ˾��x�&�e�����D�,�<����㨀;"{���L������`V.P[��q$.��������b)O��;6�4�E��d�H���#�+JyY��!��ǃ�2*�Ѽ�ƾnͮh�F�tKRR�Q[��	�"�ZM���4����� �j'�C��6�Xz��r.jdb-Q�_�Q���-W;W�����Ҵ�ۥ�T&��w5�1*p�ˌ2���FX�NBذU4~bg���))	���:��tF��.0"�������$2f*�0�!�a�&�3i�nk:8��3�3�����-�9P��l�����lN0D�_�}
:����h���H�H�����`2?���)�x �*p~�Ml��b�=a�bդ�.��-͑�����W�z\l�R������s'�����̺��X�����\vg#ac�/�b�G��I��4!#������5�m�!!�r�0F��kI��2^�:FM˯����7���A�8�iu���ŏTb/y���=�l����{T0Uϸ������/�1�a�ۯ75C~o��B�<WhH(}�*'Ǟ?���i8����`��*�f�i���^����zS����s��`FL~��'��%��Kc۵�� K�(�W�}�bdJ���� 0�&�F���BjPL$}H,Ok��n�x��.�!@���T)�Zӳ�`gkS�v{�]ee��nu������-)�N���Ŏ��e�=*���Hq�<YE�1�5;���s/�:����0�Ӹ��r�]3�(��i�c��.��k�� @���rlP�۟�Ow�p&�E��L������p��mr��:��G�+Ǽ���:C|���"������S����r|����z*����-ҋ�v�s
�Q&�_�D��̉����4Ѷx�'}�\?PX�h�̠�Ɯ�?�BC>����pծ�4�i?���zE'Wq��5�Ba*ތu�#"����T 0���2��e�g.�!��J��֝���ǁ��BaNK�xX���d���g�z__����+���IX�4��T\T��7�4&qs��8S�8��d��19~r�T5��wp��¤Fv8�\����Ϛ^�l����6j8ڞ�X����U��׋I�@�����gh�܎��)��'��kS(��R��?�JlSYH6ea����5���S�eLy����͗\�y0�\J	�:󢺬�*��b��(>i���/�
��"�|���j�0�#�9�/�F��J� Y� �HQ[������Ş��21'l?��ϴ �s��~G�;N�&�@�O�=�"�y3��Ӯf�e<c���Ɵ�a�޹����s$Z }�`Ц(����fC2���XԴ<PDS��A��;2j��dl���G_k�	�lڿ<��A��l�i�����Ȥ;C�����/f�c�4��.})"u�pG�W(?.p!�
A����1��O|
��F�^�oI/h�.�֤�: �' �����d)/���3[����+�����-�1n'���ןm�&��}.��WGC� m����vܺ3f�Fsw�,���C��I��y7����%g�nvQ��P
��D��Q�ϥ¨���4�A>�A�Ğ⽏�nzzT��٩��|�	��%����s$�BI�:V���\�r�Oxx�B��j���+L`ߡ]r�.q��ڨ0z�V4�ئo����_- ��Aƴ�9�&.W2��<�'��*�8����M�].�k�ʞ�f�r�B:L!FU���9�`A,�MyN�pA��=Q���������	8Ƕ>�|qؚ����W�"�G��h�i���� љ���Y��E8_���n������؞�6�PYA�B�6ZB�H��[7��O#����7ko6/	���B#]m�D��P�.N_����f]b?�%��iM��_����U�~����*#� ��C�;�2���s.���'.������5���pM�����I�DVL���I߭�C\�����
�@~P\y�m��~��ش�Ã�T��RԂ~��)/���#k���#�߰O(�z;��K8��6�5���
qtFf>�Bs���˕-!��2���?]�L����0 ���_=p#n���A���c�ʙ�Fe������Z�ū�� c�+_.+xF��T!�Bǯ!!ͣ�_�i��������SOe?����ڳ6S���O�4��=
�_�Y%�w��	�b��8��q��S�O�̪��O������>*�̀"��V�.� ��ֵ�O���;;ъr~́Qд{U�����J��F�sD� �o��.@J�C1������j����P���T�I/���`����h�0S��,3Ǆ-�hE��Q����!� �v���)�N:�&G������ղaO]�ۄ&�=+C�����W��/W6��fL��Ca��?���%��vN�n���#KƂ/H����ہ�?{eʯ� |�x��ܯ�9<��"��l,u�t�R��Ag��\N�/k�$Mj����$m�w@�q�/���sф�~b`�X!�{��.�s�f|����z�{8��+���6��1J�o8��z�}q�#h�ſ1d��;6}��;�Ap,b�ܟ�I��󣇮BM&��[���zk)�ޏ���5q��I$k�O�������t�E�F��0.7�g Ϳ�H���?E�L�X·��`jƶ
��er���:�.:.���O���{��v�g�F+h��J�T�)>|�����r�������������q�N��P����k�p�H�E��^|��3� -�&�e���Z��&T8�㎂�P��ޗd�~ٛ��Mt��g��7[`T���_Y� 0���I��4C��uoĿ�\>��H�<ݩάj�!Z�	���� ��ĝ�$��b'�u�G|%d�d�ಂ ~�	�<7J��[-&A���œ��w�_��$����R�)�i�����,�C;q�i����=:�`�]�Ȱ�����k�\#��C�_h�t�"�v|�(�&�_ٝi�v��vh�)����jI�����]
|�-�h���I��_b�-#�N��Y����F��p�\hf�OȐ&��wc۬�5�@&�WT�~�~����0��
|�.���3���員A�U��y������Y��1����%9�-�5~�7����ɭJ�Ls?��䒂��=f7Yʩ�g�$L7H mFk�؏((:)�gt���ЗSC1�o��%Z���df�{�U0�a�ڨ	@@����3)��hn(����(�F#c�Y�Ig~�U�y\�-�Qx�VE�i��=�'��h$̲�=Q-˾tDsg����Dǫ�I"Z��=V�V�pK�|:_�9��,Z ��;i��I�`pqu^PBrL���Vc��a-�~<jp�t�b� V�ƃ��M��*���c۠�(��N�߭�T8V�p~�G�a��SY�[��tP��佼o�눆���j�H�gYL�m�2*��<�?�K��:k��M��$�7���ӭL��K��,��xU�%R�����(Y��M> ��6n��Pm�+������lq�eX�����nwӦfe�����ft�܋یsW�m���|���X�{Nu0���d3����
[���d\�D:�o�lfSp�Q�����ιZ"s�=U�����NL�݄� .~���$�7�eC�3l4˂���dj�@!<��u��r�����o-�Ƣ�S<����p��;�;���ؿ' �7�C�� ��E(��q���\�"S�>�s ����?��9���K����8�"hKZǵ}Gu~MG@�'y�~c$+��]��)��a[#������
d����1��>]�jH���X�|:�P仁Y��Ul�nuehkiߥ�/�����3�?�2m�0�ߚ��1�8<Ɋ"|+���p�=m:'
y��~��*�'T.����Q{�y��BoѸ3�Vv�qgr|�-߁���2�̓Ia��yޖ:j��rc�6��[z���Ȣ����[�c܄{������h�q�഼uaVU�����:0�z��IN^�����X!p�"���d'� q�?N���F�����&��ge;n��O��oѲ:�~3>�O7ˠ����V�\�@a�|�Z���AQ�o��_���ino�&��Kh3��e|�Nl���͕~��C��?��A�L�D߇�t��CeY����O���*��y �x ��̞� �ݶw6�T7�����s��b?+_��7&ɐ���5ċT�����f���M�6V�T�����]@dݣ�8nև�f�\/��� @�#S� u���V5�۞��
e�7bS�z�x��*���r�d�\��h+��$K�g�Eb�Zgq�ټ�y���['4`S,����Q�#3�(٧����Z.�0���E���)K��9��fD>����u2����^� h㆖:(�)3s��=�B���#�$���m8Sxr���Ζ ��}}l�R-t�G��$��4��޿��L�Kv��ïB_?�0�����ڀ;����_�:�'P����J��(Ec��ư:��r�sq{��ɠ��������|����_�E?�~��]a��n��R��hL��|NbU'� vT,к���/)ps �3�������Fe���sP�T��-����e�g5�f�&��հ�/�.uۇcI��0C���h�L�xZ�`'}�uą�p�jr��Y�?0h��;�|)0[ṋ�:�ģ�K�Xk�|g��E���B��N��{%����T����DEʼ[�R����@�!f)�a
���bD �Y�K��䞨��쀜��5x�2�p.9U��[dج�Iv����&#L��ϕY��9�L� 3,Zҍ��Y�X��K�����t��v#�'�;��+���4p�Y�?�� x���V2�&wS�m#]J��iH{bh+�w��4��\۵J�j�Q�SS��L�37�n��;���[�>��w�lN���Q&ҁ���g�V�^�g��ܣ��v��u}@�%�b�Ph&(�	�)�cHM\'bS�E0������\T~����񆻽�b���MzGbj�m���e�k���z��yO�m5JPu\m������0L-��p8�A蟼��R��tS\��-p���m���� �.������iY�]v�����b�FH�Gn��(7k*�ǘ���Fp�*����F]eܪ��3K�/��1�i�7]����L�������_�镢DM��v��L64����llnq0�Q��gK�$&����As�� \W�;]T��� ���R����g���^��q$q���m��e�s`gF�-.}��]jVra���ƺJ9$��𽌥#n>n��~`�v�К�`�e!-ѿEA4�I�x�+������Tb�& ���-��΍��l�Sf` Y)�ҩ�y$��E�eo@���1,����@G��}�@<N�?㨃�gv�6ا£I���s���&�������ּ{[�$g0>�:YLD=��-qAVD`g���c��<Z,lמ�gK�5Z7��1�YX�xe���nxB�#' :�O�����#��E_%���ͭ�a�i#�ܬ��A�8�w�͐�/#4����������ոZ<�;>,�Z=?�{!0�b�I���,
mNE<[�T��U{�H�O��<����5� ��"�s�z��վVԦ#1:�@\5���ѣ�a_*�3!�G^RXd���Y����]�c�/u�b�B\bQC�\��>�4����g���}��S�o0#����8.+��R|��!I��X�l�O�3�|�*��Նr�;�t�����Y��!n�C��w��=�E��$�XN�����
_-�9�� ,T�q�ܴ�y�ӂR��@��d��X�z1v4�}	}X/�r�l�tb�F��M%-�͒/�$wv&g�&��p#�����n*>�%��x����:r��=�����K��ݣ�LaO���j
���Tp+�[MD(�\��#�^x�̓��z��5�SԖZ�����s���b@�'/t��;����f�e�V�o@x�nҬ�"Udw[ �h0�={��V��|>�1M��lVe�����R�"%��tv\Ӹ���2�K��tw2�Z ��fC�.C�T���{�s�QD�f(�o�13˨�QTZ�7K�{��-����t��(�|	{Ȍkt|�����0��t3��D��
8�=[Ǎՠ�k�E֮3</¿� ��=�ϰWV�х�[ˡ��i�/x��ܬ.=k��
��	�e����Cz�9���a�1� ht�]�BN��Rv)$v�v��������E�?���~
��i-�H�����ph����q�3��
�.��m�N$+�d�/ ?ℍ�������&p���R�<�� J� h�Y	w@n��n�E���'�)�_�J�W"�GP�T_�.�Xj��8m��p�#�f��O��"(���ֱ�I��)vA��� ���k�0����ʱ[s~ŨNj��Q�@{�݂>P���S\٪��W�NLIS'���*r�g�6��W�Y���3T�C�����	�öT������L��p�ũA���v�+Q*YT�r#[���)$���ߗ��ݤe��`�����(�n� �C���ت�bNn%��)������ge�,�m�rt���`[TY+r�a��ܩ��Э�����g-{��Zj��I���WT����h���Й����U[�'�Q[����b��Օ���3/�7����߲�СI��,�NB�R^g��� K�g���5�q��9�&��S`E֒����m��o�\"����6��o�h�Z�(J�&HY,�\�f	~2II M����jo��WW0�?ǚ9@\�[&S�_����Y�X�9��9�9�n��T�2�/ϙ>
�M��Ϗ��863�Hv�F&��4p�gɯ��r��4:$��˝�d�Hf�N;����_�����u�M�/���K"�Q��bQs n��q�1��%��t�߀�@@�$�Ր��DG��o�5V\V�-�} �p��\�C\v����9���R��zK(:��~J��)*7Q���7���M:{�d�/L�7�Wۗ#g�5<�����n���aD�#`�&�"9�=抧0(SP���y��K�c(2�D�y��<��c�W#߉���ǹ+rx���>�����s��-�� Гx�'�ߔ�ǝ�1P<T�WH04?��I#���?b��R]ב���\+�K+&�F���ǀ ��^���_�����Ԟ~�鯇��݁���6�G����&;d���
���n9�v�I�����v��{ޜ��v	�&��`~q��3���[���ei/��y6b��N�kW��
ޭ�"J^߯VF�]�x��q�$"&��X�O���(H0�9l�]�;��� �?�9�SU;��榨�<d��(O6�1~`��i�
�M(G� ��r^�9k ������q2^��H�>�"�r�`����z��,��% s�	�����{�aNp�����L�PP�-)���`�i����$�Þtr}>{lo�kŴ^S����PΒaڀ[��.���' ���z�-V ݦ�g�>Eѯ�Q$R%���dj�q~z���]&�!nsH��=�Y�n<Z���M��G����1�B���=�Y�U/���&�A�.�H��w5�K�($��N;n�g(8��]���A�9,�At4���V��}j��؅覰n�+م���F�m�_���*/����sf&�꺢� �j���eZ��|z&�	x�
/�R��4LBN*��a׃��y�/$� ��j��R��3���)�>�(�=���e�,R��ZPŹ���G�o
��g_��6s���	ß�d��g�����	n��W��}5�A~{��-ƭ�<X\��w�� �}TW�5>ܿ�����R��@_�����h�&��@/f!zyv�Uwa2�o��t����D���F�ǃ�1]7��B�ҿ�>ߓ(gu0Ͽ|�!xunzӘ���f�b�,oW�m�G��x�oN��������ycR|E����|3뭆�n�E<ίa�]%�(��F��p��.�{�4�Uq!�>,R�)k�����1ǟB�jْʹ[�n����x�������A����`k�6��o&^���ʷ����e'�-�t�U�(�F��7�~���d���t��^�9<���'����s������	gcx�4�a	�q@��
������<���B��*e�7���B1�A��_N���=�~��P,r}ciK��	��:UKd�#�cx(��C��}�Tܙ{1	C���A�d����ƀ�j�j?�pt��g6'�>�J�5�.g�JPb̯HޜW%3�����c3��[#ˢ
/7�Q�cP_t��[�(3������6X�O�7b����>Z��]J��禺��9��>��؆��#����#�D�"�z�>�����e�?�!�����[3��2鬃A#��=|�����˨
�� L���5�gi����=,l���e\������NH|�k~�p-�$/H&f�@X�{���̡Zt�%!�x�G�}+ �W� ]�D��a٫װgǕ�RT��v?�!x�*Oby4A��&����9"�l#��� *."fg8���ih��
����t���1��J��bt�j���Y~�s�$����n����X<�8~�|Y8)�BC7�à2z�!�3A��d���Kh�(lz�h�����{#�W��u�h�ƫ���q�!0���6Tv�!���Ց,����B��=ܯL��U���j��zc^�2�f���I�m���B͚��>�k��5V��XH���8��3���WȒ#툊v6�ב����>n֒��yf��AX��o��,�?+p�������:"��?�Fw-}�-Dl��듩u�eX_��8c;�~�T�߃&,�w����l
�q��HQm��ͫ�E����z;�_�iCM�y��6
C#���@�^Y��}VdV(��a���zLr��4����2��ZV@�!�,��w
-w�;�"�,\ɷ7@������	A��oGf�ik��k6	��;j.x�a��)�U�K�98ۦG���kGp"D��"6�p�ی^ni�:��!&E6�~��O"6�'��X>X��cLȄK�' �۬��-X^ l�K��T�e��<�h�^��M3+���0�Z��ag��*���tb}��Tȩ����e��u� �^�^����'����K��ɰ%.��ٛ�z�@^���MV�%�:��]}�#��S��fb�a� y!�N�o�!�9������·xl.���vÌT����$9�i��5�p�l��u9~W�"%W7{ �Ϩb��"�&ӕ��c�՜S3�&�x��N�H:�#zIڅ����9by�݀%�0=� ���朊�:�%�/Q�3ܐ`Jo�y�ΩN ���nP�;yIS���<�����v�KI:"�2jvEi�9A�{���=3
�Nz����:�2�|���jvi��+�����T���j<���|��D�!�b8
��b�VS!��i,,J6N����1������3P�2%0��,���{A�M(vG���^��I�����z@��W��\o���AY@�j9���&������y�Z�k{sr��X,�BV֮�E�Azl`z��z���a���v�1D*�r��d'��:�m*�p��z7� Գ�rX�z�\^����BPY��aY�9
	�|�G')��G�=��x���iPuDЈ;=,��ﯟ�I�f�|G����Ma�9b:��@
m� �re��$�����6�a�/gD5���j>>�#���a��N��$�w��(�NȚ�Csj�f_Z�㽇\���;�cg@�џDDs�;��*�V��x� ���?9JJ4��4�X[�ycp2�'����9�?�'����g�
��/l�9}HUQ����1_VE8d�^�e˃����s$Gw�_�0�SO)�0d����Q���7,O3ɍ�K�<�a�Z��qǣ�#0[3��7X�b㔦��Hd��D�e7pc�ŤDJ*�'�rMT�����b ���A�PIN>��Q�義\8���?�e��z1e����m<<���&�m� $�q��#�}��D�N��M�S�� #��|�؇IRm���k�ו�&�w��IzM�W���8|�oG,�g���w-z��bGZJ��c�D��x�U��ir������jڑ�ћ�_�D}0���!����1|�K�O��D�6�Y�,O��Qz���}$ؿ��7�6���~4�.!q���j<V4�����I����/�>`2��*` ���{66�5�7�{�s�A��(�����Bl�-'�.�@J��ވ���-�i>�.�g��ڵ��Æ�0�G�W+�ӥ�~�|U;��K	n�/���H�Y�O8�F�?؇��	�LK��{'� �\kp��v*�����*%⡒q���-��Z�xOV�j
R��A�e�8����z@z���no��Hv��$�3�������g��맬u\�G1l!�=V\c��T
ɘC��Gyn�< �p�B�<o/��ɘ�s{��C����|��1��*gwO�?���R1~���r[���X# ���h��j��V&f��;`�$q�����s�������\�<k�s5+Q_y� �nG$���M	�Lg�P��NJ��R��>��N^]hi�H�8h�:�v�7�1��ϔ]��{teŲ�*e���m��S�o~�t��O*��!]����[�����6Y��=	��-Z��]t
�E�8X�p*�$q�y��ft���W�Ząh�uH:��S���B��$��梽�c���	'[�Y�ƌ����"���r���i8�񢢳����[|�V���s���P�H�)#�D���������&��^W�εo����>?K��S�UR��&B ��z�����CW����Q˺*�x��	4��ޛ���Q��Ϧ�w�o$A5��p�'���Y^폍�ͱG���(~��V������jް2~���%���2���@��hbH�
�q��w�_�:���@�o����س��M��z����WI��pz<d��v����[�	ᶳ���5�Ӧ�+$���u�g�i���=�p2b����d� u�V��Wo3'�P��~�>�#5|G���i�J��Mt	GF���w�D@>�R~��%BJQ2.ݨ{��'L(�m]Q[+���v���*�����C��^,/`0W�&�L��6�ؙ�-Y���9�h�(���{}�,˪ȅ��| 	4X���V�w�^f�Rn��A
�y˻��B*?=f~ݮ�
�~��x�ȓ����̋�#Im-�p�/`$�@��R��da��7�$���J�qz(��ɇ�XР��k�	1���;G��M������^v�4���E�����{�	�}��6�����2���fQ��5��j�l��&�<�MZ�DG~�ű�b롚�b�}�R4`+��(\A�N`�C��T�:���\2wt؃#7�f�F6VV����ک�)�J<��2:pN�Z]�]��t�8�$,�WOu���c�u�}�>=�oCd�Z��QȮ�/��ꊬ�`���pM�/���ᔎʉ�	ۦ�(I�kJ���^��Щk�g7�\*d
����ceO�W� �(^��ӰU�/�����B� a�0�J�6C/0c��f�v\M��xivGh��l	��ɱ��5��!.ٮd�֧6\J��W���u}�賩2G��.ҹ]^8,Pf�m�J�y�U5�J��T��Ap��k�����ܗ�
���x��4M0}p	2��=����K4`�ś�kS�yeB���J�V% V��B�L:��2LN9�Z�r��.��ԇ=�`S^qA�F����tsZ�� �w���2�#ݚ����7ކ��ޣJ�6J�V�^I7/���0�^l쀊��˹0������?M�s��$��|E@��|.M&��H
�]
�;&ݶ��^��َ�\���술�M��H�����$�?4�M7��@���<ϼT |�F�=�f�՛M]��֔I� �����s�%JN��JG��cֆ��6��	��-?��
�D��\�h��S��b��Aq��pb��X8�z�̗�"Z3z#����L�!����^[��':��7�d5~�;I��z��Bj��(���$�;���[t˙�Ɇs�k��0���e�P�=	SN��[m��K��� �k��"�0Xe5��؀M��0�l�5���G�:�9��Л!n���`ۧ8;��K9@�yd1��9:NdY�x!t�w�KJ3��P���H��y��?/��88Ò}Gd
�U+�CNt,�HՂ��&�J��\�i����AN����a�1/�p.�2q��uC2�FdCڰ�-Cg}$i�.8�>6��#�g��y���˼oWg�/H 8�$�QWWGr�����@���ľx��A�p�QV)��_�=�~��iک�b8����x��2�������-(7�>�(�S�[ɠRd:Rв�v�����Fq��k^�?Zl�s�	��4&�Y��&KU�QR5.V�*zb�S�����	���-��k�?�f�۸�ưu����t��u/�(ܣx?o�ӑw�����xA�q���I�e�ɦ�Zed����ՐB�pԃ���Şw�ct�[��%.�ݴ�c�Du����ixh���N�i�׻b��(�'la�d���;
DT�sC����Y�t M.�䅧�ZiU|���nWCd��f|M�d�P}� ��,^�]ζ����g�T��.
�Y�����@4
�A�A�FcI�����=��p������:��=-�yD���0 [W���,�rw+�}�@7���G��J�W�="-��?���O��O{Y�~r�Ga�M�9�H$g&�FLg�=�����C��X�P�؝��K
�3�@JGOZ|#W�d̉��H�)�
5bX��I]p [F�p����7x�:��M��J��s�H�}�\X�m���	¿�7�^�����4]�y�f��|�Jd9��k�1�1|�fjql�Yȼ��PB}�R���yE���5<%Ѩ��"�GNb/�����.��(�î��E4���u�y�0H���J�F
I��lf{VC�ñ	��8c8�q)�ҫ
="�K�r�f��7@��J�c��憧��!%�y9kgF3]��]Xn-����M�l,5=� t��&C�B��)��_���	�@�(�QH���8Z�X\f6,=��iW���l
��K#;���'�c����]K-�e�[��:�����ғ�k�˗q�]��w�^����»�p���*���7	��p�@�o%bɔ,xa|�-WZTl����~���]9�Om�dR�2��H�����:Z�4��
�-�#�乚��z�H�� ��Ͻ�c���+����;��Yv�1�F���MvvK�,w#JMk�\k�������v��chG7-���rH�묗1׭����3�+T�t?$��BV�o2��aRu�>��	����]���R�8�,��!�?��j��k~ s�в�.�s�DhovVHS��󂹶i��P����N:9}�@`�|&(Ά��
n!�(��0�4�f�Zt.b�u�o!�Jʪ`�U�R�?p���p�hM��Q�vlSj}��&}�0�b��)�����ȄR-O�G\��MiF�8M���]��w�v]RNgU6:Y�ܦ���雊1�>�j�om�#����/2E����(�QcsL�1Ə8O�Au7*��(�����kqx�K%}�� z嵇\"�m�J�7��´0��t]��Nj�O��C�8sW�.�b�}��9�t��_d&�RL��:��P���;�sl� 8ڋ}g�l�#���'����'�����a�V���v���j����y(Z.����>�Z��a���+~CNi��@�FVH��о+S*�f3�l���Q�����N��Ȟ�3�����ƹ���fI��-��$:�Z�"7����)�۫�J���:/�]׻gm�ik4�2GΊ��=���>�a�`��M������k���َ��4~��5_� ��	����(!?�Al�wWp%Ҵ�.Q�3l��y�0f���!���sպ�_Quܵ
��JE�G4̜?�aY��:�gʩJ�x�'�wݒ$�.�Z��ã�#{G�U��X�+A�%��Gy�Q[���/Llf$V�%�HX�G��)�-Q�/����g�u����~����D4N]1Lk�8c���q������tI�����Exh�c%zB��ۣ����a��8�������Sf�iKh����s��Cm9��%ޮIV���_�����9Q_�84��'Ҟ�Y�T#�p��wh1ţ|�Cy�Y���(ny׶�N+����x��jX��*���tgU�$��#Mi��� ��5�?B���}q=C+��N�ݡ9��_��g��߽�Ô�'Q�'HZ�v
)�������M�i0�R-��3%������ьiP*;�����<��I$mg >�q'�0�Tc�t(��2����q�h�殻�ȦM�F���9l����8�=��߼�BB*F}Q����|z;Ȭg�7g$l�c_��h�,I,A�1��(#wfU�]�	)|JpT���%YO|�[�����y�k���%�%�4�dn]�"���by�DU���>�|RYul��}X�c!9]��8@E�J˹�b[�;r�.a&?�g��-:\熐�i
z_��X����������1�p4�^��Z%>5���� uT�꧗�'��	c#��ͨl�%��~�s^�Aڌ���"�i��<�l�~|,��r�
�jE�;&�����}�Rn�l�{|ӄ����A@�ٜ�G.=�+%������4�
���T��Mp���y'e�'ĭ�P["+m`~���=1����2^~z7r�#OUM��[�V��Oɕ9ez6�g��zذ=o�5��3H�\O9�q���]1"������{Cο��#L��&4�-f�~�C&'Ջ�N��g������FOr��M�$Ut-�qT��/z2Ldn��4B�Z;��^8\Ƀ8R3?��.�Ɠ��HE\BejH���`��ؒ�g�:3�ѺL^B1���^�[��^@竐��+�,M��L�o��ν�W��A xGs������)��`&�]���}�/;t0-����=1��=[��}��o7�F�3_���d����b��!��F�+z�u�bV��ͫ~M�����_ZN�鱨$J"�Ň�ҸKfm9�o�#G�M������	�������9�E��\�ǌV6sј����a����"��Z��S��t�^�Y*�|DԱ����v�l)w%:u����؂X�\���BU�Z�n�(���n�m ����R-i2��̙��8�9X��ɓ�N��L���T1zlL��Ү������{��Uo�Zq��*<�xf4XSBS����$"`Z��� M�S�J-��:�˿��d,�
��V>�8��Ҷ��
4�E6�� Z㩩1i9���B9>�[a$�6F;(��I`�,&�J9XQ��9�vRZE��b���Krb�D��m��������7�̒�K�0j�{3)I�'q6���v6�R�ڡ�2\�����m����(�r���+M%�L�������w��nN�5riS�Ws/$b����u/Xd�.��g�
���$�M7�v��aCT��c�G2�s>�C;}@� ���0�A"�;�k�|�������9?�������
�MR�\��χ���@��;��c� Ϋ�o^|�[�Y����,���e�ė����u��KK�S��5+�Q*&���=7�O�-U�*O.m��L��ቁ�+Է�O�묍�>�p��5�y����g���~�ۢ�ڭ������E.h����k���&vl3z m	]0��.4� �RrO�c[��=�~g^�c��0K"T��-^�,]�˺��z>K�<EN��6�:�Z�f�����ji��B�
�+W��-r����O��(f�5z��Ȏ��g<�Ux�܃/#-��*0+����c��2qg�B>�C�"��C�|��}Dn��&�#��S�{��Ʉ Jc��&�"-��#�n�w��5
�\�����d��L�-�2��`�+�k�9��E+>O=���9��빏=����_����P�Z��DVu㉁̓���>�1"�i��/~���h`��"�H�d��A'sA�j:<睱��R���W�����V�_b��ۥRe6L�W��3p���c�N�(OSc��oՠ�W6����f��8��3e.��y-7T�b ����ǵ�-P�sb��Bb���c|Ǧ=R��MpA�]�'�����i��ۃ�<��|(�y6�%�,���SH9����^;X{2h3�=[6��h�GmJ��z}Q��_Qݏ�]��NW���^:��@tɁ�9�y. ϠiT�r�(5�3��j���5���#�rS��-2���.�D�����or��]=���d�sVEk���u���]�Ɠ��6RW�'iW�F���^G|�k�8]w/��ŕ��)(�G�G��%�T��$���!�,�rsc�r��Ϳ8�!�+�=`4ES�j����A�[)z�7iX�����vuC��r���A.��jp�o���˽G	�H4��-}V�B1mӾ��l���E�(2\�>�����c�k��٫S�4'��V��h�j��޲j�ۼ�3� ��/y�[o��m{mݥ|�S �@�uC@�W�tlz/\�޶rK��ͯ�o�k�p�Ð���f�me3�p�и�f�!�y��}��A�x��
�a�}: B#��wv94��y`�)�c���P!n��,��uhF�aE���b���9"���X��lN�ɵ��9�Hr:ץ�(jz1a�*�9�6&�o�`?��]S�2E�d�,ۃ �=Ê���Qj����l�6����Ư\�s^\�-+ C.Q�;գc"g$��7�1�X�Y_��q��׬BJ�����KA�/�uk_�g�G�GpG�w��@ L����1�܃���§���GND(鶠����H3<��6�_-���GД���W	�4c�c`�9��c����o���&h���� ��`���me{��wq�yV�>�ѵ��7����۟;}�5�j���u�D��f)���yY�s���ʔR���^%�'δ�տx���vz��%�|��EWpL$���5kf�{|��m#�xZv����kBw5���~�^U���b��ˬ���^\*	�?wќ�dyK�P�5B�IF^%�q�|}r&ԯc� w���nt�����P龅2X�[�c�~�^D���{	���>�e��g]��*0��Ņ$x (eMC��F$B�zu��f��qj@y�0.��4F���v�২t��L�Y�?w�����m}xpF��x�v�M�<z`*���H��E��?�r�|�-�Ad�(܎!K�!��'o�����S]~,
;G:����D�`"��N��YO�1��c�"�?;i�B5yD��b���r�d�9Q]4Oa��|���YY��;���u��s��ޏVh���ƾ鱿yV�_q1�E�͏E�,��6>���`�������iW8�h�?>�IAt���4w��GP�+����t��x����-A�D\���y�&�Ь�#o�0��2�ٹ��i���h�c������B��>a��ͨt�ir���n�L�G
y+�i�5��Ae�\��N�� ׺���:e?��˹��rA��vΑ�y����q먍�r�Q`�(����d'���P�����`&��b���#����܂�n������H�톧O�|=*�S����3V�3 F�=��V����-�5
K�~Ld�k��!|a#\B��-˥ɋ�l}��ě��{j`���.B���8������p0	�-ޞFU7�a0��I��ё.^Z����-$���=�x%�Y�_u
�3��O�J�.zA�8��&�xGWAn�+�C_�[�"3Y��c�+a�߃�3	�ě5Z}r�Q�X�������P*��V��F1�˟���o�7�/�Iw��9�\��;���8��:n�j$'��ǜ��檣���F�b�*?����/-O||�p`R��4?s�!����{1���D��$�����6
_'�3'���#I���V,��_��5�1�am�)�-��̈�H@K���a�Ei�d#��\jFv΄]~�įDy��̣��ֶ�������M\U!��MN&8�,
� �>��A�T�?����D}�V��є!���Dy���J�Z������ZR�o��#�N-�
���^�­&~<?�Z[P)���
�;Vbpel�����l���K�^�nF���0���÷��J�2�����
�v�M,b����
ᖡ=��HF�����㓱Ԯ�|w���A�ʕS	�0|Q霹� ORƜ��kw��{y��l8��+^��˼u^!�& ����ܪ�x~�߸�S��,�����">Ύ���3�l���*T�%d��ʃt�֮f<���}�9�w��=�L1����'ֶFG���0��v$�\�a�0���Ɉ�$z\���!!�z	�y?�.M���j���3�u��a�z8�ۆ�L�_�"��"	;�?>%��[�a^E��س�G1K�[��4"��Z����Ɓ�e��ݼ��O-�-���<h�@�O0}�@�]��C���c����"&Y�לi Ar���x��O��{�ͣ ����7��F+��_{cnH<�I`�^l?H}��hv[�huъ�2ۖ�r�~_��7|(�a�D:���B2v�0drȤ�q���E���}3�H�E�ƞ��.��Me���`]���s-X��[�S� ׮��;�4�կ�ςC�V�Ò�0t��,�?$��+�4�|�[�=9�:�tFS�A�m��|�L���Y �~<p�u�s,�i)v��>]n��+kzY��Ia,�(G��C�6����^�`�_	Yf/�������b��>���<�r�T�DF�C�T��'U�/ʫ ��c�{�F���g�����xݿ��ǰ�����Ci^�4�'�������x�_��4�H_\� Rc�S f��aO�N�]Z�RX�'�����ci�]��P����w��h`�Y�?����C��	0n+���m�y	E����&WvvS[���v4LӜb䈐��Ľ��sgʎ���.�|p�?���/pxn�]�x�w?![���{Gzy�:�lg
Ŕ��T�!�qr�Y��{�0r�O�T���(�������4Qk)��t
�-">����AC^�����ݝ��(O��ׅbE[�۾B4��z�ٞ~�#t)������4�y�����Kq"�	[�}o����a!� �}ۨj^�L�IT��a��@���$tb�[��>6r3��ަ4EaiF���v�\��i�́�n�f�`���Ls�<=]�*��Z'�ri?/B��$E��5�,�q=^w�HP(��,�x;^���'����Ox�К��*PP���9^�H�w�{Փ<�����=s7F`m?�0���2�!a9+�r	|��]���"󧻵�����̪��
��߾�L�C�A#'���5-X�����yp�_5�p��	wŦ�\�9��0���w�`ɖ�<�Z�oA�4�K�XT�U�U����F�����^u%��Fǉ� �Fn�by�!����&"�P������m��
飚��9AMhO66�0�w�,r4U���G���ӳvʩ~��u;;s����F��e�����Pc����e�/�c˶���yb���[so=*��Ձ$?��`��}~�!X���������=�HT-/k�����Ʌa����Q<�����E����l������i9��ۜ"��d��;�6���Ä�u\nc�w���p��5�4���[i��j>E�jJ�NZ�
����u��*����d<@�cT iy��E� �����\�/@�/�'�ͯ��~�F�'�zG�$��0N�fH�":Jaٶ,��g�vh�O�9�>y_-B:v4��դr:q=�Q��BHv�5�.{.-��_�o���n���HBpC��|���:���� ����C���3����C�;H)�D���1�1�J�S��ki��r�p��́�����kda:FħU��uڹ���0��"�Iz)�ǃL���YjL��s՛&4��
Mzb�2L�i���M�E2O��C"��Q��n�F0<��v畖�a(��`���$��&ɠ��*�*Q�N~��=�ᣦ\Aj9އ������~2����'ǫI)����f%��5E�D���l�n��
V֭B����50��$�mr��#;��VґA��7};����!��`
�~��F9���㩲�N�{�]�\.RJ{.|A��7�G�X����m�¸�]�ppFX�C@x376ڤޭ���\C���}����Zv�"d��``}	��+l�n/5��\*�I��O��"NF�u'm�3���9/�v����և?���kd�GT�AG圊M�1]�t�h����8
�<��.l�O�Z��B����̘<o��t	�v��[獏�T�{L��+#�u�����/L�9��8ՠ��4�8�h���Ks��`>�Ԅ�0�	χ�Cp��s� g�>�xޯ��o��nrDc��."J�N4O����0bO�LǣT�H�>���9N��	����0����7Z�)�G��p��	<D�ô�;��?����������]*7�TkYN �
r5�xƛq�TC��ν^���Q<��"�l�;(��� �DL���/6�׼����>�u�1M"FRAG�8H�<�4�F̰R&"-��&��"EmdYY�u��N��@���,{0U&�=oň�x(/��D���.oŅo���	� �@�sTs
#���� "��q<�$��
�`���+FTA�nȝK�L}�n6��p����Q��D1}Ε��s1���^���l'�_ݡpb��H�s��+��� ����+��r��F$,���O�')�F�1��A%?����]�<};>��T͊h�O+{b'��N˼�7�=����r��K��5(��$�h��s3k���/�c8|�Lx�;���R�bus�	��BEhѢ`͚������K�l�0���.�(;ތ����շ��w7�l��12I�H�Vy����� r\�@��{����[�%@6��"2���z~�m��].Ȣs�e|��	��C��Ǩ
)y��Qq�!�cٹ��v�J��S�/�	��u��TW��@(�Z� t=�X~5�c�tAǐ��!�P�o�'㓗6!#��ë�:� �H����	�Q��L�5���^9���5�Q����N���'A�A�F�麴��d��uz���H@C��7G�
�YOdi��Q���P�� ���,}SLA�N7��v�f�x�j�C5��8z׽�~5/�0�����9�Te~]<.{6��ZЙԦ��"�O�C����9B7��;��%���O큤�L��{�}(a53G�/�5#W!+�j�͹�����ln�?��lb�ѹ�]�;��Q%����b�����{�f.6%GJ�6y��8]N�}Qu�}��v������d�����Ē�I *�d>Z|y'�P�/1�Bb�|J��C5@�&�+Q��צ�rs��1���F��/~�[�4+"����+��<������#��X�� XuQI���Z�[&7R��r�IǉÍ�?�h����;��8p��=��C\�Mc�m.�~A����p�M�����p�9�R�[Y�'yϋ��.�����
��X�������T@�=�Bؤ>e�2u�}y���8��-�ț��)�|y�tߪn#�;�@̷zA��sz#vK)����>kC�6�E5��8�5y�1��PA�U�T(y:�vK�KTi��gz�t����Q�4���}E�y���@��1Ў�[�����2و�1v=�̃���"�&%��US��V��K�ٓ��r�s�q�s������֬��9�N�c��;E��7�	^F�w�v,6�<�u山�z�bWl�����5CX��*���~��Y,I^� +�TZ���ǠRm|�[��Y]tT�����������(�5�F�&����џ�<̣.�L�%>pB��ӋP��ro�9��$�	2ZO��G} ��l< ���������Q��rl�p�<�B&�%F�Z����P����x)}^��mʖටơ�1Č:�3�z��\�F�؇��zI"0 q?�rt��ڝ�3#Z�l�=�}�ҩ�JT���	��/�'�A����ʹ{��I��OL� ����wS�1X��F�2R���ع+x�C�L5��"���p��@F��d���3��q'lL���(�Dfy��3�����P�(�A�!��G���^�V�sˏ��\���,P�z}ïIe�d��~	�p$?���♟�ӱ�������y��Ju1`,Mp|�!��yۭZ���i�6d���5U��#�ms>c��'q-~ �_�64Ie�����ū8�]���]g���ij8d�z�>"��
��;o�;�F�ps1t�}2�aZW�8����ՋR#V����:1����M�p��=FP6��X��xdeJ
���"H/KGB�ه�3)�7�J��ы�8+�)��kM��ۨ-����ϟ��lӌ&MG=+K�*�e�2qJ;j!����̺z0�ۃ����5C��c	���i�mHK3�f�sW3}S�
p�?0�6~6������E�J		�{u���%ڻM�5���Ԃto�H0�3�f4	sI�:,~�1�T������D�Yn���27w�Ggd���E�w]����V��)f��_�>��w���-���l]�c�p�_,h�&|	ΣAsR�w�~�u��X�����o}���e�.�N>ޱXm\l�p_�wCt�i#b��Ec��T��@�U�0+���$�jzry�S'Vi���`qy�f����
�k�����w��h�E���`.��
DPV۝8	�c��wa�!��Wa*�����.�����F���Uk�y$�{9̮���\����B�oG*�Smh	܆ �t� N�5D=}�a�r��QO��f�&��3 �C�K�)�Ļ)�KKi@muSq闻 �|8y�*��G*��ԇ�	�@
�׭7��yax@ۺ"��w���oc;HGl�BJ�t5@���{N����c�'�q}0���*���S[A���*���V�B�����z�8�ߝ_���N��@'4L����m˂�}S]��<�i���b�h�6B���U���E�:E�U��3�m2
:O��s�����M�5�R�^Q|G,d�WQ����bC��nז�J��*ޕ���c������?8k�ƀa?얫�J=fX�+�(��M��M�,7��)�zBN2M��j�0�ƍ"~�q��:I��G���N�K'�S�T�n��F<�`xZ��AXݜ��J\�C�ѿLq�ʋJ��%�MPx�)��|o��T[Ȉ��TQ
�;��QU�V��Ml^����_^��1*"�۲��}����O=x0]�q����3���ʈ	��MxJZBރJ�D�����`g�ٽ�3"�=�e٧ �\f�a ����_���νf�k���C�=��D�)!ٶ2�a����j�6�ټ�Ǖ�鬝�������в�������9?H�]�ȵ�0oQ��7�O= i�x:4b�F�s���`F���0�+5:�Z����(�{��	E���8��e��2b���_Y�<�����DX�}p��+�d�׷a8aM�T�5߁S`0=ZL�)���=R�n�t٘])���t!�ms��� 0�l!�3:u�}t`���Tgc�t��E�|!Y�G�[�Qu˫�N�͊B;��u��c}{�OWL�X���kR���j�B��_�(}��m#��nAC��׼S4g�s#'n���$6*v
����"hP��EZ&��.cE���ʘ��4���A��]�)ͧV�A��N'Ӳ@"������;p��Yc2�dZ�3�ⲽ�O�H1�7���W�l6f�lĵP%@�����C�4�_��`��B�?��s�����\�f���������@_
:��b�X(qp ��PR�_n�ګ�qy�bk��%�����p"VZ�ڻy���Djx��&�-7��[uC��ϣ�eE1A&u�j��	q�����V�캸��
l˓�x1���1d������Pzbc]'m��G�~�v��F�+$���RӔs��P�)鲢|U�zd�)��S%^�2i���~8�<R2%5ǌ�����i �v["t0����cu97�TjԹB�����=�AV7�TX��M���|�
��7��ǎ�#i�g�0^��A��E�P�*-;��2��>7\���V�Ժ��HUF܈f}��4&�����M�ȅ�c T����岬8$`�&���{����Ut��njD�@�W̍;t��t�XI�R��)�;i�\���r7��͙:�Ȇ�@C|l��I�ٍ]S�,�����Gf-�Г����8~�5c�-��p�Hd���V?�LO��dN)�*o��gi9���]$P;l��H�;���ط�/*�+=í.KW*l���R����08G[���8�?��+�����Ɣ�w�'aYYVTs�?�y��9�y9ѝ*�e��-�8� )5Y�K����.dS{G%ȃ� MH���6/���&=��RDo�R��z(1&�ۜ�}߭�؜"�\~Z���r�
��peկOR4����NI�y�Y���!�������dk�ѵm8���4�����wŬWQ���^��z$!��徼%�BД�v����s�$�����	�5���Ԏ}���-`�@���FrB��Ƽ���U��f=�P�4=��]؂ӯ?q��7�X�T�0b�Х7(�a<�U	��������w FS�2��ޭ"[D�^�eA�ߜP���D��z/�.�=yd�}����68M$5S��k����s1��0�ĉ�2Ym�i)f��.<�����ꀸ�u�b,h�q�iS=���	�Mkf��[PI&�NAj����)ȀY�]��E`L�{������m�&�c>�����hb��<�~FQv0'����H^���cu�]���c�,_�S����b+��-���(	��eb߀!�Xߥ�����ֽ���Oy8T�e@3�m TTbY2�:ȘJ9C�����%n�~��x��
>�/�&b���W)�\%I�.r( a:f^��	s��y�M�[)7Il�"��_��l�^Or����-��5�6�ɲ9hC�Q��I������U�h�Z��T0YO~'�#�%�3�7ލ���{�Ti1P��]��MD9H0F��֎���IE�������]g��Ten3�͐!�1�~�����Ӯ�����s�̹�hs�}K~u�Iɑ+�Gj�O��F�8Ц'. |����n�!{��e��4��MYTv\�k{�FR��1�b5�P�Q�z��s�yk�<�$��{wE�6�GY���^��_���~]�����d�u���GZ~�����ђ��U$��2��B�����q�z�I_���F)��͉]øY�K\�~|
��KmC=�0)�Q&�ih3��P�2�X��JH<VK��������~xBX�'�0E
T믿BVU�"�i
�fߵ������ss%�~��q�}�B�p�{e�iZ�srh|��+��2J�}�Rw���F�}��U3�(�94�����VL��}	�$^��nNA?�G�1k��EC�4Q��<�3%����Y�G�� e ��5ݞ�C����;S����)��(��%�Ut�L>Q�R��֕��i+2���$��J�ߕ1+TO�����$u��,j��c]
/h����s;���J�	a�.
u�u���-r���N���� ��}���� ȁ�c�H�q����u՛�&���FlXEVry�1�SgJ�F��B����Ԥ�$�%XbF�H�!�p��Li�C��,h�H j���ݾ\�~Gk�g]��!%Ҹ�P�ˌh����� -��Ϯri53+�aD��
i8.�06g�����S�0�Cv>K��	
U�k����)��.}�p��N0�5�##���C ����I�fj�=��(F��4�X쪫�r�М(�l��w��W�]�Ub-�q|�E�x#
�8'C@��t}� ���p�Y�FM��D�'�-�yjY�ɬ h_���ޙJ�6�S�.\V���4_"g<e�U��M����f��oNc����f�|.�����(�xu�v�<���H��n��윖�bLx��v_{?�(U��{���ƾ4V���ݗ� �Jog�T��!��)���'�8�<��nu�0���.����Δ��tל��R�w�R ����e6�{�(��C�@Зhu��e�Bٵ�[8�|zD�N*u���g{����J���as������șj�!��w@΄�T�*�K��a�p6X�f��"n�~�?�=d/�~2��[s�V��g*��w& ,�#G��-V���&�������֭N.K��T�Ds{�W��z"�?��-Ϲr��5ϧ��f�+JsB2����Su����;\^TY`E6xa��:N�$�}�1���J������,��'�o���4`"�{;C����kR�Ye,;����*v`�u؍@��4Z���G��$*�כr|$Q�kx��`��:J�@��^��ne�Y�2Ƭ��,ˢ����H!�t�6�� G�v�E�$٪�����<��'x�gb��JI�ڴ]nw�~���$Gf'](iW��']��OT_҆V�,q榏�$G�,�8]gJ%�4�K�8dj��`3�[2F�f�j���_�z���F��@Y'�l�g�G*���$6i;��%�W����X���:���~*��07�����v2�ַJ�f��t�/W�?�PDF��r�u7D
��R�ݵ��\]�U<���~{��
���O�N���=,�R���;⨢n]5���l	���Q>�`��^^@���--X&�<���{���������6�|�N0��g2Bqk�r�t�6oS���^23���0����/(+�:ϊ��(�"����Y�|?@l�aTj����L3�Xg۴7݅���۶2�_>��B+_t�&$R�gT'��VEp������L Q�V+�'��B"�̳V2B����tT�koh���	�G$S2��^���'�:�]��fb���#����
�֕Y��D���2�4��`?[�F�gt����X���RO��A�ޥ��`�y&�˺
��լ�2{@ }��P@�|"om��/_��oD�R���_�t������#�΀̏���@PѲu�VT�1�e�� ��I���3�u�иT�#�1F�$�%߇��?�a�X6��Ѐ�p��c��3�"��i�+5Y��k���H�+�	HC/?����u���/�y70�d��5���
�B�:�|{���;�B�K�(e�"�0v�σ$ q�BT3P��E�[�ـnA��NP�PT�m$^�R���.lu-{�`���l�1���;`�/�̷!�Pgʈy�7�^����B���P
Y�i�b�I�\F��Ϊ�fYؕ.�&�X7�!R|�.��$��^V�4�b֟���P�����4F��3���}�!59��/t�Xj��m��J��Q��\<��%�<|2RbR���7̻.�W���LR3�!�![0ɕ�r�Č����V�q�7�MF�zB4�W��n��ə̺�<F�I'_r�J���(�$����k�g�y��3D����-�:v���:ChP�TF���ü���"[�xӏ񰰖c��I�Y��5V��TË��6���;9 �l�x��ڎc�<�Fl�9��8��h���(1��tl63���Y@:�ïojHR>�#����]L��j��f�,�;��
�/M�R�G�u��a`6$*%��>B�QV(��v*C��KG9Y�;�mƏ(�/:V�t��P"ǹ�ԩ�ּ���,��g]D}�m"� PXQoVV�u>h%؜���$hu4!�\ӅTP�.²k��B7B�;#H)դ��Ó1q!sϠ�����nIGQL�hpx��i��VN��U�,�fh��Ӕ[�0
s�����׽/G'���:U�L�:e=K	]�6�c_���8�K*��(�<�V�iX7 ���s8f�>=��A��<61�?	�DS1o��a%�C��������V੐�#>R4�(� *Ut��о
\V8#��]����)�0���>��}�U$mJ��1-�Ș=�ىx(�W�ӽ,�p�D�X�E��0��Ғ|8o�0g��!�p;&A�L���i=��9�ʜ�W�f�3=*���5�W����G��M���? ^�7�$�[_�Jen6R� �{Pw��qE���NX������U|�n����߲�3�WOAnq�ɡE�Rv[Xn��䥗��j� ���|�>Xa�6tH	9��u����z�`�4�.q��Mc��@(�8�^E8G�����k7�CE�ϣ�F�m�. �9ґ����UƝk��:=�:u���U=۝�ưF�Qխp�9��K+l2��2�ATv���-��2j�7��Vn�'�t2[r�>��d��!pE������z���͞��\c�AK�N��0a�6�����{����S~���J� �y�]�u�z�Bj9���,�T��P}#���D���fd�%��dd�?�{�6RaЖ�Q(�X���K�']�@׭�Z~I��ZF|�Q������+7�o e�g-��Uv\<^� ����K�`���Q���6`����w�V�k�����7����٪,�=[F��)z�4��5�C$g���� )�|vKq�� �i&C��t�N�G�?��Fׄ���ۍ�b���=�	�v��I��u��r`�Ӭ�����D�߁�(� ���֢q������wOg�`�ccN\���ȽS�A��jB����?��~��ɤs�%�I�̰�EE[፥��p#�&���6�?[�Jɼ#��R�ug@$�������Jg���$�r�'�Ux��]$�r��K��٤#��m��=c&$ ^�bi�R��������%c����K�k,�����{ʢD�Jy��3@$t6sqA3��5�w%���<�A��'?h@ �����Z��L�%�v���)��q��)Uz�	&_�?�a#RC���"�������i����8p�.�Y�-J�vN�V�y�0ףbFS��aP/���1ir��;��Au�v��f�/�9�O���j}'�I�?B�G���j�߈�~�D-�Y<��<q4��-)G���BX�j�_�` N]��`�}#�!��		�j��	�Mh�_C5gF����2U�wi���ٴ�o��P�5%���3�y��?�?/�k��g����Z�7޵��[L@+�byW/��d��|���l��0�,��a����iT
��k�$PT���n�����S3^�aؤm��J����|�b����r}S�`��/�G&�UII�w����J������Co��>��b$�O.�G�K�롎�ba
�g>�x,��@��ݷ��X(��.�\Z�_:��\��L9���w���T��.K���.p��C'���E!/f�=���˓��[�:�����1���ZOy�0�[k�P?	R�E�P�j@6�#�q5�64M6��8[v��ŝf*b0,��Pm�w0�C�2��t�k�ȑ�8��@�����F�z
�������
Z��;-��y�Ӵ�[T�J�s���S�[E���mV�w�؃��#�~�`;�S�ItYDJ<���w���UP��򥊯S��;��{E1f����V��:?��1ԩ|0��2�oq��W)}�x)��Q��_��� ���C�$�0����ʹk���˕�(��*�CP�FW��|ϗ��ڕ5w���
� �ݐ��u�[Ya���qy�j�s��Fd.*J��"y�N<��P6�/7���p�ֳc���>n
�"������#�j�wfJ4�6;1�`z^	Mj��s��gA��L	<^_��l�z������y�@&�J��������ov����jV���ޯ���hz��k _U�E�b�	�ݫ�h�ax5��A�c����ˉ��J�r;�Qa�ʰ^@�l�H�6�Qh��Rd=�G}��:���q�+�4�����Z9$3Ir��|z��,�G��N�4�S<Ǽ��t��n�����'{���ZY���'3�|D��i5J��!_�quӬ�v�kH6���L���O`r�e�b�=���!&l���?�W��S� 'Kׁ�	�X�Ə�h}�a6��f2s�lU{W28�q�R�_������'5 j����É�~]���~��*%�4C�3�W��EHHGa^4ts���S��s�g>�S�KV��Ev�����2)jK��r��h����&?�LQ�BC,D�B�S�""�0p�RH�QH���+eOX���4��)�D5����j�I�9N�Y�
ϋ��r��^��ΐ(-�D>A#�Ba�րi�kb��5d�Z���͜2���8q���S1d[�5�u#VY�z�Cׯ�B.����3V���`��H4��x7*���C|��Ǫǀ
�r��(hS�T����:C��yf-;(t���X�{�lܻ�O>���24�jp����ѫ�j�?�9>���c�z� gq�����<Z�)~:2�ǵQ�j�@+_�s׉�H\r� ]o���+�ƫ�T����^�z�����X/���&�y��gxWh�L$���M�nR��x@B��L�8
��Ǿ�I.π�I}��O�0�-g��s�o8
�*��$�w>�����<t��Y3�i�,_h����q��\X�է�}�����bK!O��L��9.A<-Mx�����׀o�d�����o�3;Y�!��qÙhY�a ƛ��Ӛ����v�_W+mhV�3�]�����$״L����E�;��hM��ܱ�?����D`z�'��N#���	
D�/���,�$�����%�,M��4	]�ܴ�3h�=3ŭr3�ץ�z7b7��bٞ����kP�[�b\y�2��;�����r�@�
8��6�����ǎ�Q�+½���c����L�9��K���=����\m��@�l���em�&�T��!���G8 ����1x��v��sz"�w��=*dK���~Q��r��M��9|�t�2G�������R�Y+ɓ}=4�0o��̼���NZI�`�r��P�t��z�ypڒOU±�r�A	W��Va	�h!`�Vb9�>��#�#м����e�Ȼ5_��%�@�J����L����Xr��x�[��T:p@7���(P��31��؃�Bܧ��f1TF�T��5�f���n�������~J^Ps�/���8�q��1ÊEH%�~�Z��zt���ƿZzR�>�=q*K�O��_����J[�A��{���M'����^K,�'E2�i�`�Chd��WDΰ���|G�.8�9��?o�*Ru�<�v�y�������`�)�"/1���k��@A�-Ӎ�@��̳�*�ș��f��8�N��R��R �Og�-F��
�����}��к�^4���Ǩs���j�S� \4��q彐�GpW�]��d2�'�5�����m��9t#�\ӳgl��JY%���?�C<�
��IA]�����.2�&
u5�z�G��f�G�����8pP,f�w�Pp�^���������jӔ�}��1�C�dՙ�/�W�)�$�5o]vυ�a{l��DΖX�r�JCr|7=S��E�T�vH.��(>8&>�geL��S��J=-����7��銡Q��d�X������_�[Ls��]��c|��¸/�u�Wzf�;W�)�#��* K������`	f]��6�׆�4�&:�`UOT�T�z��C<Hɒ.�@�I$��`����$a$�A��˖v�H� �W�aݒ�<*���Ƈ2&;(`�����]K��lJ��z_[�6!˚TWWE�V�yG�d��<�۩{xm�	
`�V�l�{��j$��E�.�Z.���� ���_�=�%�i�	7j[Zƶ�B2VW!#��E'L�<�gӾ��Rz��g�<�	bc�v�^��bK��v���:7+$t���}`���2����a2dm�� ��ׯl���D<1�0�1�=���,*�y`�]P�ø ����V5��n���U\!*1��'R��5�/#(�i�A׭ɇ@�l5����&�~	�V��$�6�Lp�h������M�9+�" m�M���MzB�f����� �RBdW7��^t��+��h0�`� +�c�*������[�Bo�jYn߉�b�f)��F:��ߦ�^x{��4;V��7m�j��,�B9I�I�ЃZ:��2�� ����2#'��m��cg���jן�FԦ�H����d4P��ݝ]8�-�YRW�#(q�ϟ������TG���cXd� !(�ػ�۴��D[�νыf[H����?���`�h���YtB��1ߢ��$P�oܶ�n�,5q4�Hb�M��?�](T;����U��[4]��W}|E�Z�8���Tv�>=(�ő�/�`�{b��n�vސelÃ��T�e��,k�@�D�k�����E	ǲL�(\�P��C�G�<��}�Δ,MojB5�|�XҴ���96�w.(yO0ELMa��u��a��k��j$�p?=�ƈ��*9�;ܻP+l����8�N���y7�'�&�+�6|��a���=�y�/3���:�*����L��`�n��	��l�1S�F�|�CEac�\DjRz{|�RI��^Q���/���d��}�F
c��AKV˂rÿ��L�4��?��^4�:&N_-^B�rX1ގD�{T�6�tF������$�&k��|fU��x�T �6���x}���^Oim�$.���"�d5�/�e�l'��B8b�N�����=R��C��ߊ#M��0�/K�$���PR���]7��BΚw�J^�'�G����	~P��K�����j�,0h\V�Y`CZ}wV�	BqǢOie(@�ɨ'�]�2��$q-_��N�7��H�f���G<���O݌'@C���n:|7yy;�чۜ}q^[��Oe�ǒfR��Ȅ��P%AF�@�Bo������{�n��3�S���h�_F�Ckl��Ҩ�A��]�	U���x\�H@�\��{�w`�#�
4�tL��=��O*TD��r�A�r��n�T}3�����m{$�,���>sL�<��1�5k�g�nh~��ql�sk%��Ӎ��e�E~�����%��nmŇ7�-P�2ӡ�[L�ဳ;�e���g�z�E_䕿�,e��(�n6���6�����c�.q�h �_S1����V��.����@G�N�9z������������E���%~�:��반���兓�JܓYz���AO$nl_��N�/�RC�#��=.��~��8��H6���*�pʏ}p/���B� Y�6��('o����>�9�@��w];�nK-�F1�?���>G;MOn���1z���
C��8!�����-q���X�"D��x$���&'Q�O��ž>K5�P�{s�G�D�<UII��I&:�d����qPC�����gLp�(���$l�(̞���뚰q�y�cƙ�Z��~�E�k9��
q�4	��9��U���q̾��ZCQe|�l�_D��=�0d��۝X��(�s��C���Ŏ����6ԺzZL�w�'�* G��)�bO�E�f��y����w
z�3�F�i�ڗ�ygA��$�^�Dņ�󴌾Q�X�]��Tر2���=(�_RY9o��q�x��9��`��L��b�����W�1���&���Hqb�?јmw�>>#�KX� �qu��2�@�_+Ү񑑚;����3��߶7ּ�
���\r|s=ecm��|X�+�6%���	P%1C}-诱$�2=��3���|�Dn����`�v7�n NKH�s���/�߆/ڢ�)ul7f�C��|L@Ld�}^kf8^��oG�Z0�(�hUNޣ|Vv~&��k����c#udQ�`�K.gS̻2Tz|3��7S��61��C̕�;�!}��҉�8�P��&=hC��D����!��Z�}Dj!�.�+}����1�x��ta\߫��ʛ#tֽ�rԪ�d�"[�F��V�u���0�)R�� |і#���Uq��؍6�&W[V�9�Ĳd$�B�N�N�m�KyD/v��&��/�OH����?wv�e�9�(ƩJ	��J\u���eG�
uKk��eI&������g�֒�x�f��W��t�H�� o� ���(*��S��}?��~�Pt�~��נ��57 x^��u�ܨV΃�&�!FV�dɕRK0�@�6� ��I���/�u S�_�V[|����,	:��&�K������Q�U��s!�^�(8����l�S!*�8`H����W�0�_�l��T`����J���z�W?>��d����r.-���_$FY~ۣsKgz��D���d�R���}1��JT�KW������YY��ؓ.�"Tї�'��s��+@m}�6���W6��p��KȨ����m��f�K�(���rϘ���8��n9�B/~����C��j��� �D-�s����x�����L��6�٨�u�i�������ULj�(6��\��ޜ0i��Ju_��B�Sl(�ϕw�U�H��[xl������P�+��+��>#�߁�nC���@�S��,��8�]i@�A�ko��£S��.�b�뇦�c��'y=M��п��]��!�h{�3���yEj1�H!>��k���^�{�O��i�SZI��ߟ�������t]@U���	]�2�t��,��ÀʗS]� �����U�8���v��U�/��W�9����ggLD٦�/'�|�SZ���� &#�D-W� ����&]0A�5�TC ���?�Z�62RR ���&Dtb���A��.�נ���4���@���m ��|��`���8E��ۜ�{���/���t���S�ʈ�`O���ĥ�0���Yy3��,&t��t @��U?�%��ۋ�x	�-U��p�w,a��kVl�X Y�Wg/��C�ŗ#��5*Ɍ���C���]6�/��R��@.��w�(����D_�j�j���R>�R��ًQB�_�v;4��S�R�&\GU�_ײ���KdMI
i������Kv�����إ�q�S�&�5�4�Dy�rN��d��i	L��*�����r���}\��X�0���A3#^�'��u4�����ow䜭Tʭuc�6�B�B�!~�Ǿ�;W{��uk!7�=y
~�)1RM�tP�9F�͑��k����ӛ�?��Gnŷu��Q�6�W��V�`?��|�P4iH��-�8���**��h���o��)��E�?�g�[�a��R]$���"E���������S��D�a���ćɱ�T*��ʵ52�ᒰ�g]nf�y'�b���"����l�n<=��d*��F��_��|�n޷�	7F�W�&�L�	�vXD�&�}J�5Ix�!�0X����pX�r�D��l�������;�,td�Rf����}���o��98c[S���I�O[X��D3|#`�M�	Q� ǒ�����o�t�i����: 8�/8�"Ğ���>0���o ݧ�bm�_j��w�F��A�q�"�9��x���ꗬ�dSu�������1����5�ml���wβaV�S�؃��=1To�t+7U�7��t�����a�����*.��%y�L��y��8��p̓j�Q�S�\g�$�l��Xr����"���{�z]�4z�<��ܿ�`�������V��K��M�]�j�4mn�v�
����Ց�Wr��$�A�{���]�
����9I����k绔;�'WK�0����h�N�xUAa���;�=�c�����ܷNI=����[mS(�?l��!`�̐�Y�{�o�!�����g���o����o���d���U	-kؔ�Bt��H�ǁ���X�`Ij���zo�m�Ff�R�b�O/P�c��%�9��;�m�'�ɞ�h�̼3)��R�i{��i�łތ���XQ�}s��/�p�nH����/ �X���C��ʱ�)I��Z�%�Q;���
��J�Ǩ�8y_�g��������M��^�|x5���������MO�����n�°kw�2�q/��Sw�AZ����Av(ǻCIL��ȣ|�ّYZ(���X���鑭��K�:ű.��*�/v��4R�A�$�?����h�q�::j��*X|�G��7���LOoeƗ��p�Z�����@Z�b������I��
������f{��f<��t���E%�w@�N?[:�^Q\9%�����#s�Y����-%d:��'�Y]Ɋ������	�K:����>���a����\�3��P��U�N~��.�����#���iK0���Cu�ŧN��A�/e�(n����.�!\f%�����}��@ׯ��=�؏H�j��5D��x�|r�)Ķ�}n8����|h�CVbH�g���t́{��+Uގ�ĠB��H�
�n�/(p�B�Ǒ ��$
k�彫�UV�k4"V�RK�m�a����H9K�����o;o ���}�?8��mN�'|���������-���� ��ԼD�����Q�h{Y@v4�8H3N���L�Spx�T��G��~�� q��\;�.Z���Z%��#�8k�$q�8�(��&k H�Y�sY���ܞ����臐��Tku��g�ĳ&�ci���B_  _U���� ]���t�Iү ���>@v�l����0[%��{`�*��Q�U�������e�# ���'U��(܅�ԘK�4� �������[���
�^�2�`-�x�kH0�3�xj���}���o�)�gSh[�*F����I��sfow=�tƵo���6���v-=�s�0|D(�h�*=wو���,�����D^U�S�C}��5A��P�` ^ၘ_LUJ�c���F��\ ���ą�D$�{v�L��X!�e�N�߬Haʢ�X�	F�Kg�'"��Ҩ@v�~�ZpF���T2�����7x�I͜W��j����U�~�3{餱G���ݮw���R)l�����Ù���C;
��Y���(�&f�^Q�]�[l[���L�.7_����P|�׸�
-�K4����.2�Zѩ���@�W������C7(�f�}#�u��E�_NG��ҫ_gH�:)�Z�e���o�C�]ּռ�[��Øi�y�G�A!E,����?D|*��]��B�] �|�sҚ�{P��1߲'�na@�"	������p8�uG�QpC�����Z~�����Ŕ>�\�����F�jn���q�>0ufc�݃"\�V�������<	j���X�"#.�8�	�O_����	�=q�W]�(&l���I����mi�<���9`�a*Y�s��)(��cG� �4��܀�o�B}y.T��$�=�gXo�)i��Ҡ �[  ry�� @���;���Ѩ���i�s� �a �K�BuDo�x�,�󥴛m� 2��bG�n��3�Y ��Pٺj��[�.�L���橡B�K�Y��|<�,����Э s�-д"��jVs(
����i�xbK�[�H��B-��=�;E��s[�S�uW���;}�6|-*p|�_�+/�!���X�a��f���Q���)xp�\ٴ%>!�J/��kp݈��}-�7F)L_�i�G?���xr�^iEf��C+6�P���J�� T�?!�V�f}Ʒ�tmBť�¹+�+�o�������^��N4a��gT�\�;!WP�L]=��Q��wv+���`KҒQK�:: ?Y�T"�N�5�pܷzi�o&#{Xj9�"$ݝ�ST%�y���8�y0�њ,>=��y�Ȥ����4�`О�쾂��y?�ye畤?�jF����7 �WF�Gh�UF��+ �����h���pR9lY%D�AK<��>������B��?��+�M8bI��r�]�1���� o��07�dgz[�LH�V��N�D3m}�R��r�/]Jn�*kҋ��qZr�w`4|%M?�lpc.�h"W�����H��,��&������M�X���v�Z���bq�z���kٓ�A�7�`--XM'�͈D�X(ؚ��[�wL�f: �SH ț����!��N������g �P���Ga#h��ǝՌ�%&�E�:r�l|eK�}%�yj�t��0P�q�70�[���dc�=/2��mFC~�%;�Ĵ��MQ�w@�a%sq��d��d�YME��v��1�`A���3�:i�Aw�iWɀȼ��V��>(�*�zN��Li�y��עv��;�S��a������,K@�!|���}��k���+h��@���J�����d�^�!p��]���{�Ӽ�b4]��Ut@+�#x��h ��,�V���פů����+ 8��~F%�w���K�<�r$�;�(?]�R�Y�ձnnq�M��_e�id���S?z��Ե`��=���M�gv�0�ϐvFV��`���:�ԯ͞�R�a� �e�1h���Ǖ��%��q� &����r�F&1�'��'�����p;� ����.�T�#����Bv����=]�fh̪��<�Re�"#�QLP��V"�qW�L����g��f��,x�~ms7*�Ȕ�Zs__-[�_���O��0��ΑD��4������9�]Y�V�>�)tO��Wa�ߠe��,�hϴ����*ػ���`�K3v^��C�T��*p w���܁�PxZ��&�{�窹��^�	�^����a��{`L�8��5q���|�������Y�x!2"��e-V:����İ�yHH#9�Uf�����v�,�c����k�-�(I�1I^>}���l��;�S?ڸS����4
����_4����{���K��C����%��/�r�iŁչ��h��Q�í��4 ���F��N`�Gi�Y�ڱK| (ZU)䧘L�w���7ƈz��T|
�L��2]��m��.}���x���'�R���]�Jx�4#9�S"�&e	e����N�o�l�ݻ������'�}
&G5���Vq��Ь�s�]"D#{'�Xz��lh����d�w� [+�FG]X{
y���<��$3Q����h͋�BWs���'��+��W��=b#���ˇ=u<�?d96��Y�;L�N`�r��H
%���0c'v��J�%������\��X�ԑ��l�6%����sD�{,�^�p9��(qY;H�r��S���*��߅ꕨ?�U�� j����y�a���c�xM2͕vBf��VOBm���Q��!�\g��u����cE�{qQ�kA@S��>����l�0���Խ{A1,k���V��͍���'��>Vt��Tik�OY����2�YXK���E��H��Qn��-�!�B�kl����BH����HYBX62�O~r����n1��B��]jޯ%���8d6c����0`�,Ž�a�����5qtS1 d.�TvӨW�1fR5DF}ۻ;��;;�f���s���l(׹�|�t��ɋ"o'yw���%"��ה;��̰J;��f^��_�Zh�X���r��=���x���5W�^9Pʐ a��kW�fRo09/C
$�Z�e<��`�N�l5a�r�\J���ȷ�/��`���5������I�z&xʷF�c)��,z� ���4N�.�����\
$@�.M%f*����9Xj���,pptC�Gd�6�F�"�����p������jZt**A��w�( ��@��B��.z~��ƻ��ز��3E#�h�L�ܕ�(Y{iL8��)��2\���W��u�@��;2�ڼ�ҏ�B���)��J���"K�1�^Y��DJ���:C�C,ә�1UR���%��C���`P�>�X�ƃi�����7d���y�!�KJV���gs
>V�`�'4�VzRa7��i��I���%NE�`�����V@ѣzT'�cl��0�6i��o�N�w+�q1dZ��a�Q	Hu Pe��l����v�fލ��lǶ};�^CbÍ�q��Jѳ�J�o���eQ��g���4�0-�ܫ�_\�K���_��n����4A<�C酳�83�A�Ϻ�1</ At'��P��!��a����N%�p4j���-�?;��7X:�,�e/��)�r|R�s�|�C�w	6*8h�hR=Ď�O���ee6|ig�ZI=\�Ī��!-��v\�l�Z%.H�&*�c�l�>��&�|)Z��{�� c]��lL1���O�7ƽeX4-ɳ$҃*nl�.�.�5���23
E{a����H`|;�����j��u��$K��n;��8"�oT,���L�2��)���Kt�c����w��㷰n�'Q j��k�J��x� f��R��Q���Q���j��<&߄�8`�x�i$�7�t�bØ��b�x�y�����y�~�ќ<=���<��ѩ�F���9���S��Mԫ����u�M^�Y/7�����l�@��ڗ���n���U;>����-Z:26\��ͻ�ӑ�A 5����������qNS?+�]�`�ͱ��������{�3A�0�t[���{� ]�_������Rj��E��b��D��a�!�q���,��Lt��|��V��ԞG���W�*~%�ӟ��!f�a�6�����פc@M���ޛ�t��j:}#��}��:�^/6��t��jy�.�ߙ2�V2��'y/o����,n��_�ހ9R��Ab���%��Ŝs��Zm�l�@�&D�N���p3F��c��bw<�=#��޸�����-�>� ����eS�߄u����2���\a�E���Cv꿊��P���LsW�ɝ���[������zO�z1ѳ�{���4���/)eFc��b����rg����VA!A]k��I­��zp0�=}
�O��72�y�7i�L��#��fC!;�4���t�810���TC��q�)N'@d�<q�U<E����bْ2S<���"g��%أ�����۳�rKK�Em�>�c��`��,��1��Y$%���v��W�Hc짳�]�k�k�K��F�[0\D��ߟ�/*)N�~��L!���/���R�/!��C�=���u���0��4�>��e�w�����������A �P#����y��=�آ`�$p�wK��ˤ�G�j�k�Qeg�rgD�J�w�:AK��\��Нi�������{��+vrOӪ[g�M3!6[�ω�u?��
.�0MYt���;c1������b<0���ަ�&c��`�3ݬ��	bÞ4�*<cP��bM1�s.5ɆBZ�Y/P����Zy`�*s/��0��!��f�9[Rض��� ��_�u��>��T���R�ϯ#ֻ�D%5�!�/g��?3%�1��}Ϸ�+BK��#��|(댚S^X�\�)D�*��6l�������Z��6Zj�!�p5�<�X�<AkZ�<�5��5n�����\��o;���3��o�w�񙑪Ɓ�b�T�D�vub� ���t�\Ρ;	pT��nBJ�4� ,��w�Z��r�����<��=2g�5S:�Q=�h�{+ΪO��p�7�h���G dF�1��ZE��m�ϐ�ϴ9H���(����f�\2}���|4�������b2ta�$#�r _�[��c��+� �~~�6���I��<	����:\Ymѭ�g��ö��q�:�'ۇ����ʻ1���U�p�?�8S�N���zqi�躵]JA�b9w>�i�W�s��>j�Ҁ��^�"�P=��؄��Z�>%d����7�{]��Q�u��&���\ן(�'RBsܓ��a�uL38d����@Ґ�#����L:0v�R�1�����: <&���V3�3u�%)MA�4��@F�4�Kl!c�^K�d�Ԗ�T1;�)��8u���]>,���8��LD¨��n�q�2�&��^�:=�O��<t�&[�U:Av� ����u���̱��RYݐf�
�9	P\yT�Qs���}'U�,�E��C�̰��xG�{E�{����7lK����^{�S��Ox^�����u�o;�D���g1������[����E��=��p_�۰��C��z8Z�J\Qz�~�\C/�Nk|i����˘���s.;���]O�������o�L�e����^"����Z�*���v@��N��CR��?$���{o"ॽRB��?VI�!�CrQ�Z�pEI�rA�<���o�-������}O���ӀV�TP�i�["t�iF�:whrãkb6?AЮ��^�;N\>��lx��2�1x��O5-J�����O��r5��\ ]deS�u3>�V�mW�MiM�D���gI	4��j<�#�C�ϖvXLs�[P���V2 [O��%Pj��#������4����b�ӂa5����:�y�9�3�om ������������������.�1/˚�4��0t�ۑ\�dpy@�T�Y) 3<.iD	>�	�;EDA�\G�#*�C�;��F���ij���
���e��?$=(��@h΀��ͪ�9��2}�����!��8�r���dH@ԭ阉� �X�fq�.B}�.��G�إj�zk�o�y���U�s ��Z߀ϗ����WJ��r�3�	�3rL��+銑mPƉ�3�ԃ���u(�������"5C`G�To� �=Bi��L�&b�֟ص�>�����>LS[װ��i��$�v�J��2^�ډ��Uo�P�#�����5�_1߅B����1	Ǟ�΋���T!��*K������5�b0cp��m(����k�60���1����9%�G˪8�<#BA�~5}�Ӹ�r��_.��қ�%�^�awc�|�s���Tf��.��>[�zr���4�eD��\F����ԍ��5��w��WR��D�5�g��l�UG��#�z�m�������Q-S�(V��徏C:�^3�V����-K�3?L�b�5�=S�l+��E��z��������ӹ��+P��P�[���e?�7�v��4Pi���x(�7:��А��u�>enN[)�E������]�C��O�ۍ���x����`[�i�v.�j�'��d�� .�|�4�WZL��X@��%�V�B��	xG��7�07�z{�=��oŝ����`|H<F�������_>��?�$��n��S ��`_`���X��@s��"���3���z�(�g�0����y7����CJ^O���>l����)i`�5��޲�WS'�S\��c|C}��'q`ebN�۱�P���a2�D��oQ�9>��P��-6�|N	��Dg2T��li1
���7Y<� <R-E'��+~��,��������j]�tE�0t��X�ހx�a�T5Y��¥��{�E�V$^�N��B>:	�Zw�z���Q,�5=^�7nK�jq��>��c*��\��H�y(03�CJg�h�oc�w)��a��j�2^����/��Yk?-C�B�
���V�	�o����[<g$��o���4'��#������*�s��a(N��O���z�Fd��-�(2~ҹ�X0�Ԃ�y{@t���n�������h��x��,ې�"����qv������y��
���A�� \�ۊn�f��<oK�J���T�''	�2���6�jV�S���õ�������	Z�7� ���T�^�/t\�j� "����G|C�"ۍ�c��·L��b����������vЙp:����s4�X�ɰ�<��KK��1��K]���7������
�w�Z癱8�Y��w/-���e�AW7R�S�|�:��j�G�������X�F.���#O~VYCSEO:cʢ�松8��W��c���/�ۊ�����M�!���}ߢ��~C�5"��I߼<�pg�k�>-���wO?��v����C%�["�2&�ߜÏm�灨���VZ�����Ƽ�\��UJs���C���R��o�,��1�e�x(y8AԎ��OӵJI���0
�zgp�҃�>�?��;���ymDy�D ��+4�	���d�
0�x���o7Շ�1�X�����ap�
��e���,��`�ql�� ��!�T �a	�4U8����t���#�gI1]���A�ſ*]�8���R����0䥌�0�an��^G���%~�� t���>4�eW�� �=��[��V��I�� {#�i�-���'+���F>��^ ���jT C4)J*e�_s��rUZ_y�!�zJDr�[xW��BP�H�#�^Q�@�R��}j�L�Ѝr�5ȷE�>*cNn�+�m�{Ka��@��E����}����H={�l��Q1iǟ؜�}�ʇRI���U1�B�ki�����.��8�8cNڹ}����ɥG�>�z%g�͗���"��(�֙�r�oPM�,J�A����粴x]<9Y
vh���A��6ǝ4��,��������5�Pb�{��з4�L��&y�
�SG�\M�L7�qM�J�Ԋ��E�M�mfI|�7��	i�Fq�*��`En��c��]`�xi	����Z�G.�:�	�K� ��e�xP`f5?֦�`B~�k�qpơ�E{��r�^��;¨z)���Ǒ�dūkg�����{�{��"�
~�oW����in�o���Q�)3ǘ�;�d�Zi�}Z���e��s�S�J$ۛU_ݎ��e˷���UZ5�̷pa�&�������v;�3d�l��� ��0۱Лye�%�D��Ae{�7�s@I�=�٢����@��i�	�V0u��N��#o�^T
b�޴}D���.�p�"T�qx̌-'<���}��`_\��v����s�O�$��չt���y�6���<g �90�H��H2>��LmOp��/�4���F��>e�\vD�Y�'8-�H�}g�c��^�ZgEW5�ǉ［���Nϵ��kD3�S�b�6�(���i�g�r,5�qݽ	�����y3L>�巄����վ�c�� �T�7p�'���L���w�^ăҀu+�-��i\,�fM�9y����V����5�.0��ӛ�00�kfY91��ޙW���1��'?�2��=�j�q�h���|vz�f�����
{
mI�i"�$�Op��MIP�lG�_��Y�������f{�(¦��w�PɞoNq�͈�WetV�����!�L���'��M�7�d�3&�Y�XN���j�,*�
��F�R�/�*o�͢U�'5�I3���'��k���V��Y�����%^���@0;0�'𧕬8��G�������'�^�6P��z�x���l}q��S�A�vz$�~�H$��,���\s�84�V�S��Kw��C2Ha*G���I`�8�9v��i@E(D;�v���41�=�����`<�o�'�v��LU0Sv �j�{��������ЍZ�{�Ko�{Z
v���7�(	�'<������Wo��Ē��F�1�˒*m��[y�7���7Ha3�����/�ÆT���ٙb��ϙ@��}�F��y�uVh}���oX�6	�(nޘ�t�G�sғ����W

�+Ɛ�D׸8l����~o�uW��xQ���KGM�� ?����Hy{�N�*o޶��)'V��ܚJ#<�[��K?��s���A�³$���7���g�eؔgh=��>���*��Jo����T����ݓ�IL�s��P#A)N鳦�ϔ���}��H1+!"�%���C�q�48b��C_P���f��S�c,�$(��=����E%d���A
��������A��+mG�$� ���
��'��1�1}P�z���r����R�?^]Padd�h�-Ԟ7+1B���_a��&@I�����ў�L��MZ��%�o�j�U��7�-m
g��pqOhW ΅�T@v��V� Y��C��(�&K�`:�Dߖ��O���G"�;�4�E����o��ͩ��լ��N���Ӗ��r�ƛ��S3�
��-�닚����X�ƒq�	M����ŤM5r��䫭77?�I(�d��+�HzJ�F��м7�G�� ���0[��ؕ��}��+����\!_�
+�ǻ!�P25<ٙ�Ha�C�#�i8�،Kzs}+�y��G�W�����PP��T*w�I�G�O����������"`蘍�C����ݜ����/^<��S���q�ؠ����s�>��ؿ��r�\���)�:<{s��s���Fҷ�HF����)&=:f5��p�����~*y�*?~��˙ʇwp�b�J�t4�����3�.4�����!�X��뼞�u��޶� U�ڲ�Z_��?]i��h{0�2�W�z�1H�����`�V��Go9>B����I�a�� �*����|�͎��R�����2@c��O��Zh=���wi��f[]���a`�����v�J�
�7����?�h��aEMf�Vӎ$9<��^3�'��w�Y����)v�!��+o�X���<�LE>�P[4���l�K��XefE��X0��R�d��,M��,��2��nhR����;�"n�tu� �İ4��,3  �SB�(!hiу�ں�X����wGK)%��߮�4x�^z�V��~is���F�3�����aᎩ���C�y�\�±��Ҟ�vY��V�v*s9La�R�}���(��\�;[�@g_�}�Xa����Mk3�#!�-Z��`�iQހ����vN����<�b�O��>�ɿ[k�_������cK�SS�ccJAf2�(P�3�66�8� ��0i�MW�|���j�v��M�!oc�Ј��,mv��xN�B���F��e
��/m&��5�ʫ��x��\��DJu� M9�P���x��c߂wu�%��i�!@A����&ه��?(b�2}c�t�ԥMT/E N�� �bE٣���+,τ�V��+ၒ�ZX ł9�&��ހc�jq���Y�N2Io����h�h�lP���Z���w�ga��Jn�i'÷�����&�1Kǌ5Lǭ�9g�~�QD_���)��Ȍ��Q�&���M7Ϊ���v���D��X+Y%������k%�� S��Ae��{�t�n6 R����&,�8��# ���A��Xt1�%7�7,��@l<�P�P�E�t��_� �C�^?��ԵUxK�e��k5�=^:H��>�<eB>�(d��O#nS��Z5P�����=�	�<�����U�4��6Y��@y�4��#i[y}`ۥ4#8�CH
�Wb�2�;�i��:$������D��K^�-H���Kz���^� �r4�_��M����?T}��.2����*@���1B���4:]X$-.-��\H�/kG�(�����m�	ߟ
�U��1�vO�)��u���&���6���'�ݤ¯�	���
���gT������ ݲ��W�$]�ce�+����Y�щ��B��\u��t-T�t��~C
q�&�I1�"�Ȼ��]�{v˨s;
�h�0�(��_C�+��L:�� ݅�t!采Q�l��h↍���Ck�l�!��KV(�`�3��t���H�r.C%/���&js�>����`����RF,U#zZ�Զ���"��Q!��!��:��
�ZV~D��d�5���a֚�p�}�Sk�5���$��-M��7̍�ղr���e~bɄ8�J�XL mR�[^�yA	B���VpC7?t+��c8�IW,������"�y߻9fC�A	Ȝ��A��ؗ�G(o+}�� ��c�.O��e���㍭V��Ϝ���0�9������TU9:>k�?h�Q��[W��C܊�~�T��l�Ja`T��d��'n\C-I<��cΞ?���;�O�R�+i}�U��"F\v����0�D��Ui�O��_�F����c@���EW�����Щw����W�Sy$�%�j4��̈�ݼ���=�NO'z2�tXK�v���	���)l8P9�j�H�P�<F�o/�#�����6�Wqd�re?�x���ly�Ϡ+�%�	:�����j��$*��u����&�����L"����%��e������������~y7#3E�?��<.yI�9��0�I�~��~�:����v}�{��d����p"in��,Y�Hf�7�$q܁�	2ՓT���r|��L����|�`Οu=�T�p'L�l?�8e�(�gO�U |�ՉA�&�s�;�i�����������m9�l!]�6@e����p�˩�ȴV�^[Qh��&����֘��2����Q�����xM�$�z�踬P�RHx�������\�&D�2<�����J-?�)5.�J��3���!���l��9���U��i��Z?Y!�E�
��Ant�1��Q����EY\G.�oD?s��ݦ��I��$�F�@����)��?�65�oDpx��枉���C��!ЩC΁=���ˑ�B��)�38�K3��ک>w=,),q���ϲ��A�e�y<�ꤌMD�KnxKI\��������Zy�+���k��B:}��+�<#k��&^Y�� ]a�s����&fa�I3%�x�Zd�a鍉�u�֡"_Z�EN=����l(Ys�݈����ӌf̮L�!T�� ���)$�ˁ��}��ȕ�6��F���ʅ8]f �($K�Zl芫$A��<��.��z����bTϤ��0�)�u��i�\H��!�q��F��g��p�
�f��3��ى�H�>?�Ɇ�hR�F�o�¨U���N�V �bgx��uD�WLV:�������l��)#��e-����za}<HVL_�}Lg"t��z���r���t������7����T��
gb[�3RlD�L�)J�M֊hx�g�����	U2dY�1�txv3��N�]�V��.��>@�vͨ���VE :��r���ھ,1WJg/�+����VBG@���?�B�p>�=q��&^��W���pk�~�UOT��Q�N,�l�K�Oo�� G��ҬE�����!��O=^-�X�[�O�K���s��k�`!r+
,�Z7/�7P���{
��w���[�+B���GJ=uT��-���1V����A�tt'��/v$��ג����U�K�@��u�b���Sf����	�?TGé1l^41F���MX��B�g�P����iB���q�9��%���tXo;��x��`J�Ea��|9IX��#���Xu��gT\X
S�̘��~k������|�
�;B����I��q~F���E�j��"��02�Pq�4LX��|���f���{����]}r\��5wy��2��1WOנ#�^�ǆa6q�lI���|�ɿAxz�D�c�U&]�sX[IwxZ,��SC�D�!�fu����Z�*C�'B�R��0,#�@�K,��-W�0>;����gcut��&�㯏gΒ3�*�y��m�^4�&�L��J����'���\�`lZ�łt"--'6�T��zF<�;�R��ǓU9�,Y̰2>��������p� 
��{�R�+6��b�� ���.�\�Q���Z6b��7�����P�<E���Zg�_Y}Gd^8#�I�Ȱw-�|RN�:�!��͘l��N� �ai�KY��xg�tW�(w*y�a�~������k�'XN����^�_h�嘍�`c�K�|=A����V,O���=_p��S-aIa��ݓV��)9��{[���9P�g�^j�\1|6�3����_�tdaY�`̔i��c<�,v��9�$m4,L�o���:�BPM��d�w���@���BJw�c]P�l��s�S-{�~���p0��fީ�����#(�I����%��2Wj'LO�H�AΒjC�-���<��Q3lR.f�����/�%
��,�5�
��84�'��J6��u��|X�4�����5��q4<8k�y��6�Ƭ#*!�1,!4����-?���}BPFM �nM�y�L��vG[X�_��]GGR�0�ٛ�⢶WOw�k��As�'�P	�hz���;�3Ҟ k��wI�Q����� �>��^	��_�3~�y@5Ud⋆\��E_��%"B��=�=���|o�VL���!	Yv4��9Vgo����r���¶�G�l�4�1 8&U�4Qt�?�%��	tO7��K�-�f(��Tf�ֱo����ǡ�:k%��Ā� "��!����,�c�����@�a.�f���� 醴m��v�HP�ļ0�)�����ԷQ��לJB�W'����ě������N�v9g��c���� �1P��'��}�&;̃�o�|L�k�*�����/
���Z�T\z���I�ll��?�@��Ҙ�ҥ�.ڊ:sH�V�2�c�����h���L�ہ5x�����J�R�k^X�Am����!D@�\�D�����㲴�G��*���4ͫH`�ZfSW:��>n̞��-�������7��qNY�=��d��Мd�)B�%�o_'!K��Г�i�Z����i)���'{s֦'�����.G"�x_QI�6|.O�C�H�wG�8!�Y�:��U�]�!ľ4�V�Ji`O&sڗY�V'mN�f�R�Yw������Q�/X�=�M7���+��������xXyF��+V��r��)�j������i��� ~s�VQp���G#�`��v�qC]�=���>�����2�oYq'" 6	A�����%,<D�f���sq�ٜ�m#b/�1�lB�=H��������k�?Dr�#�Z�#\MaTB��μ�`oVa��VX��#�:�RQmE���9��1�R�X�e�,�	�`���׽�1
ح�5qk���G��Z�^�����	���ſ�]�	@�(�9*^7z[r�4 �+n��Igc7=5,�S����P��JtY.�Jp��bD	�UI�o.���+s�k��p�(@IzQ��uv��%8}`iqM=M�Qn��]������v;2��#s>獀0������6���!7+Q�?��7�?�r��;t�w~�5#;v��/�X#�	 <�XG�����+�]��h�: ��LHx.i[ �Зp�8����R�!.����������;y.c�V�p��1�IZ�O�Jq4�hib
	��=
y֟�+3�<���thԿ)C2�8���z1�F�`�V��a��,�+m]E�k5�br4~���)R�0^.a�}�\R�d2q���Ѽ]�^N�А�a�
Q"����P~�#�i� �X6Bb����T:/+�dp��6���m�XS�dU�����!�pMU|�����%\���6;X� �,�?�U�G�d�+��*kP��݀_��$z��������ٞܓ�d+�Wo*u̓�"�ؗՠ�ς�0��ܿO	Dsx�Bz�����GMJ"�D��ݪP�����8��iF�_�`�z>�²wQ(��������Uw��pFK�7�+��� ґg7S|����~�����[9����|2�:��I����߱7�߆w:�G��r�71��(�^�՞��+�믱�܎z9g��cs���/Z��]�
-�%ٌ�Υ��򲤠]S�0��2��}��2��z��-�W2��I��.4����Q�?��{��U��tD0�.�K���c$��� _��וS����(0yG���B��X��t ��z�~Â�4��,꾱�$��9��a�J�l�w��ۥ<�S-R�-ɖ�5���;�!o�#�bM��/���F�͚���Йe�AekCӛ�Ql�r顗���|x���(�&�VR����7��S��#k2{b��V����f�O�,~fZ��@6����]�� �
Y�=���@�[s�U��i��+�ّF����X�hPQ�$[̈́V0D�oZ���+4:<���tq���P}I�DJ��;��tKg�h�o4�H	���f'9ʸ�O,�N{y;I�pzLQ�F�������L��9g?u�b�:���2dyR^��iLZ$,@�\��(ʤ��D�O�~;t*�di�H�}��ga_�rbD��<��R�����ݱ�
��xgD����ɂS���H�u����N[����^��U!�E2lwDc{�M>j�F9��
+�F�\���>B�7�f��wo��y_�CGb��s)�%R5���t������at�w��s�������$��,*���'B���$d�lr�C2�FцY:f��]�j�������o�( iA<7��|L�޻��t��R�����&��!��ɐ����r���:f͓e+�|�ٖ �OV~fda���3d!W���Br���#x�Z9�d�x�`S�]s���q��
AS���(	�ƭ"#��N��%��[k1ʄ���	<��Q�-�Ù��.���`	~�&h8y0OIU�"%uq�e�RY�DV�7�T`\q@6r��l����{���%����J�u���H`^��#&�7~V�J�r��$�"I��ܑ"��c؏��U3���D���J���4�^�8�����:j�OP.�����6��3_t���<�ĝ�6%n��!�(��bRS�j)�ǒ�4<�Rɪ�� ��#�."���L��x�<�O�=�(l�����1���VR��>ְ�b�\�T<��g��ƹ�w���L�-�\m�;"�(o;�\sb��T��3�cVhK�}�,G�8�g�V���t���Y��dg�`�;|
X3���z`��&��~c��z��OĆ<}�GrW�2� ��ʬ$���tA��$�~��D�uEbJ���j3Oo�m�x.��t���3�9��Å��ܑp��	8&��#���ϓP0`���v������Ñ��I�"�ـ�b�w��.,L�@_��G��NSN'�Jw5a���Qa��̠�ox��\�_�hF�G�?F8%7��Uޙ�hȄ)�",�}�fAe�`����F�S�n)��;о�C �'��:A�1SZ���?&Tkc��g��dV����n�"���*��貕ڋu_d]W��õ��{���[y�wr8�Lms]���������Ԫ��v6.�?Q�L�ptg��Y�h$����،ԉ� -���NY��Z�� ��(�˯@��1蝞p�_T5�!�w�3�Ưp�2VXC��-�-�9C��_���*a:���Q*��}`}C�#^?:NV�2�F���ƅ�ѐ�Jo�G�s�s������7�pG� #�$�XN0g����a�ep��R�H1�0g�0���{w�4i>-Xx(Uf�a�����$K'��W��*����@�CyU|�|UA��p�h�F��a�\�Kb�:�s��}mP���+Ȑ�[~�H�'�gb��z>M�N�&{/υ����l������#�Q��nn��I�����S�;*� e�L]"i(D~q�T�FB!�z� X򩄓l����.K��^��҆_��ք���D[�N��:���1��ļ��ˇ�X���rY������}�>!��w�wr׀8��Q%J ��j5��._#�(M(*I4hn���~Y�4�<�/ŵ;C����	�J�{τ�0ݓ�\ݯ|������K��vАЈ��/.���C\���C�ۦ��O	��6�2Ãɟ;���]	G|���'��Z�� ��2��3�><�Pf�:��fj`5�1 �o�B���h��d$�lJ��I  ���S��-���w�DU���v�3*T�G>8s9��%|d��~�2��t!<�;F홫�ΏA��2>�.SD�S>�nn��-;��
Ke��x7J������oQ���a�0I)��~J���Ic��j9h�� �K^�g��Cm�#)�]�V�c���9o�Eܹ��ڇ�yf`����>�5d�Bo�uH�қ� �_}W�- ��Ղ�r�9}v0y؛����i�˴,��M�Vz�H.�'�4bm)e���}�XF�=�?�{�?�
���bT�M��*��]�(H�,��Q�q,c�B΍�G�%���N�	�so��ꐶmNa��ˉ���ǟ��y���#��`z�Ŗ�~�{c�	�ӊ����Q<���S����^"73��SM���Ϗ�gD�`3)���V>��/���a%"��4��o�� ᤈ���:�~abk��r��n�|��8��	%Ke�@<U�~ ��&Ra�Zn�%C�����kR2�4��G��0 x��:����hbF��C�Ow�֙txt��4'xMrg̊So�~���'ŉo+c���Z�3��dq3�:�Qii[���;���ь�.2����u벭. �*e���$-A#'���?JȽ�����"����U<��vhG�w]�����&��q��zel/g� �uD=����zZ�/�z�@�
�3g������1��KJ���#ԓCn�,���� {��n,��K"i��ڧ�{��M��G�zko�������;=E�93~"�m�Q9w; ��T�������8'LH"�	
��i��m���h]�\�DG40"I¬a 6����x�\ �R%}O^N'֝z�g�1x�&�#\�����a�#��aZ��A�78�o���\��m�����c�ct�7i)";fW�F��G�(H�t�+WG��G|��?PY��Pxi����[���Bߎ��qciK7#|q��@�*1�x���͚زb��"E5�]0k̞4B�Dᙘ��bu̾b{�]���"@�e⅏i!Y%��ŕ�"F�*��LPu.M&�Wۮ���V�m�b�[���3G�ʭ�>�a�
�Վ#��[��"f���@�ܐ���~�j�~(桀�'&��a[�����⊙A>�ӜI�0�������	=��� O��Z�2��pS+`�<FW:��� �]>�e�C���~���������U�|��C��U�a�:~xj8Q������d-�����E���j�_�ƺ�(���U2��S��s��y嬓�X�c�	�GLX%져0c�򵁋�d ��'�v(nD(�eIڸ�i�R�Y�38W�[[p�J^i�A��,,�-�USGr��$8l��0p��M�_M�֡A��
�څ��CSq�֒�nO�Ucc �p�F���H?��`�s��oK��C�S�/��f$���KD�U&+-�5f�fi�_�"�F�Cp6l*%�>���-8H}�y`̓�6�&��d��|�G��Yns��q��21�;�:�ǄT�b9 #c	�'*f���c�`	�c�{:�MU����*�٦4D�ܠ;��4�b:ɺQ�`7~��BC����t�Ȓ25Z(z�B��9���"�e��tk�	����S%��%7�+��j
P�r�DPSpt�� ����2���5����G�2���LA���z�M��#
�jh�l�<EvX�,����g�6�T�!n�7c�^*��ag�.��dj�K����*���i����:�a\�.F���}B�iO�M	[�������,~�0[qY ���V�p ;�{6��{�p�F�8׺��}���2����gB�ϑM�M ���ޭ5������zX[uj�B�-W�2&�wu���R��ˡ��a�
7��)W}�b�E��tE�g��P�җ�Zh�+ş����ڰ�CYݮ($���d���x7S7��-n�q]p'�#(-��}K��z�~DYx���%m;�P�(�:��7����|��$�Z������	�e_��D!�|��S@Bz�F�#}�i���W���	�@�2E�UG����������A6_X1W���+���S�<9/�n-%��\Nr�\a-hvn�U@/#P�B܌Y�K0��82����Z��+%:Y��֪��`#��a��k��4l	��k9�����_�O�?�M$H95��|Uޱ���!�_XZ�8��=-���|	�j��	(���GąT<������)9���%Y#�2��?�{;���@}���(Kg��d�6D�'��S.�|1b�#/����O	0�) ����Xτ{-�`GLR����|(|� ��+�{fki�Wk�3H ��ƒR{�S&�9<���W�4�ro����Sn&��Mx��g�R<�0���oH%t�"U�I�q�`5���'�A�^��d�he
T6D��|a���$Q�!��6��4�%`���5�<Ƶ��@��ng�������a�Uk��P
�A�=�����&,A�Z��}�mD�t1X�iLr�l��\aP�8lݲH�QOq�9�0ki�5�h��_��A]y(=�9����b��ST�8��w�_%v�1�n�m�%�b?ed���W���V8�<�6y9c��nK 0f�,���9��[[R��*##Y�Z��B���X�g4#C7���	�Q�.�����x �H�N��V�ͥ���
�L�7�Z6>��{�[���"(8����ϑ4n��SXb��P�)X��l�������)?�X	�֣\�P�}'z\LNGx�ۅ;�4N"Z�=�"L9n7��K����ۋ00P�{z�����'U/����X�7*W;��i��}FhK>��'B���X3n��)BFWp�u
Rp6]�E����l͌���4U.k�.�i�j��{�W��ǔf�>z�H�Y�h1K�wF�N��ޠD"Ij����g���5��7�q���j�Tz�V�q�>�/�a�dA��RԾ=D�FU29���S�N4�U�Ef��Ƀ�,vFF���O�I6����_�ø{�מ�f_��� _��݈L��ff����êP���Pă 3�f�YԳh̼h��g?ګ�_sP��g�g��0Ii�7����~�9�F����}�;�&_��)��2�� ���P��;�5�)���bsFn�j������Q{��^V�e��� 
k�C�vHr�o�xz�O3��c����q|�^�]��,��8-���?y��Y�  ��������L ��"�A�}}������s�u��D�2rt!��n��K֗�j��>�Gd����8�`bt��\�v� ud��+M��M�y�Î��v��)��SD�ǬX�5�,$�]/Z؏�� ��N�1�F���/Mf6���۞�Z!I=\Jǟ�:e�A����Y�&�	�� w�G02���͒�m�,�X�28."*o��4{��b��L�C@�3���������7��X�k)����m���[�6Ӆ��\ �����R���]H���&� >��o�[D�J���E��v#P�4t4a�}�M)!�l{"�y63 �y��}��b�F�������I�<��f�6�sB�Mp�
ʞ��u���y~�ۢ$����΍�&BS���<zѩ�����wݣ5�OG�+]E��3���y��;�>C2�G���s�YG���ݯ�s�:�V>t����k�҉$j�
˗���Q���U�+1F�u+L�Lʵ�ЀY�'t��� �E��C��ez��Ò��6lnx�O��#���B�#X�	����A�o�u���HSFYu$T{I �-���?�SϽ�%�e����Q.�X�JI��<�K�q�<1ttf>
�t,�'�'��8��&5��2�(���r�F�e�ݨ�K+�:'�IH��.�Y��֋WH������l��!��3�^��rw�w�<o��w�3x�՚�,��;�}3"X���!Nr �n�=Z�@��4����r�����r�mW�r���C�+��k(R�-��@%��55�(�l�p���f!6?�x���d�l	'j�֣�l`�e��h<��$�l�
[�Տ)Z�����ʝ��������p1�����=�MO��=��̐ǽ�)5���dX@��ר&
2�M;�*u�扻(��I��B����7��=K,"�=*�!�j z�,^�o��J`�� گ�m4t�%���4�Q<S�
�=�t�p�I �J�EB�7j����a(��hrA������PD�x=�í�f�,���x�L<��Y_5^.������>t�.ً�*$$J��h��M�z��f�p�z�զ�["¡���٢�7��.#[�9��F�@�+rO����?���(�C��gy���v��8Yq���$��-N��>�-���8�=F)��H���iI	;h
�s��qB�@(��[�I]4GZ�ĐY�*��w;b��?�M[a��.4�h��n�9������ �#��3�b$��J��J��vcR���>�9��qGg��p�o�+H���UM���u��4�+Ŕv�:� _W��E��x�M��E�7���<A+�3{h��]�Q[Q؞��7�.'�V�J�m*P�o�R�6&Z ؍���w�q�u�Eu��>�W���r�C���]#�G&�+�
�0�=O@�A�b"���<�&;
%�ՆKl��U�ڨh����(¯EL):w��u��tؙ��;,.��K6��D]�3X"��Ɗק���W�`N��}�ȏ7B���$�Pw�Ws 8�j���Έd��ڸ�3�_�g_��)��<o]�FZ	CE���F�f��t[�����q(�G�	�"���#a�q��"E�?�Kh;<��	�|�>$'��H���cy������<Vm��'��$����J����)�I��U4��]�w$l��4#0!�+җ0�On��Q����R�lϼZ`�֘�
J��͈�	,ӈ�P�����@u	�<��ZWi�km��N��j��Qr�-)����%���N{6�i������;��KC���4��X��y���*侕pۄ�Ml���
�rS�j���K���Qz����s�ET�߭�zrl��$�-zD���sf��n=����H�_��θ��h[�l��ԝ��`����R�kF��aES�9Į�����O�3.	�P�Lޑ�E����;6���*�W07{n��p��n�A�OJd�A���=p�NUvșgY2}�q9]V�z�kҊ�5�Q/��	�Uf���V~���X�4a��]Lu��b���K���H-C��Su�*�wL%/]_E� 0�94m�����'h�Z��Kצh��TRƷc��t^J�����5��*�^�P�_�͗��p��6wn��אr_��mno�[�~��>�DV]��'x������Ʌ���3���@�P#��J\)%O������������Z�$a~��ʘ4f�+�	�*�Wa:�lXP8F�S������@����:'㫻��Z�����7�y��2B����:�� *�ӓ�'��ޱ�=���$� oA,����0{��p�btw��T���z�}���@�;Ia��2�r�E�/$�e_)F[��μ�~GU��uMXAD��"�7.��:]��~�H�#�A4�mڔ�A�%�e�a�v�҇���UfE<钾�;ZE0����ɵy�RVq�V�[��P{, u���ؓ\�
����x�F�=��Q2l�)�W�e9\�7lA��?��;�s$�9�),��$��,�<K�q�3vD��k�i7��a)"��uu`gh:���?��O�
6L��*k	�>��V��"����t޲!$1�Znw}�6�l7�K
s��v4�P�� �y�pV9?Vn�%#
rP�S����*-�L�jh����3�!��s�5ǔs>��+�8��%�c/���@��Vm�R�9���kz���^��[໗��`���-��oY����.~�_�J��Y���K++�W�G��+ �6g{�74ͣ~5����
u����뾣���k��Ž������׳97���hϋ���SM6&��͹ԫC�Ǌ����C6��R綍�$;A]�g0P��H��0I����Ƒm3���a"�7����C��-�@�	�d~��V�!v6�*즷������@a�e�������ݣ�a�-�uw��O�)�n2�"ZJ<O��\˴-H�ʦT��t=�v��M���EWt�K���ɕ��d�h�e�QՀ*%�r��8��V{�ƚ�I�_+6�.lv�SzU3���>�Ƅ!׏j���\�~�E#�f�i-z�Bj�+��-Y�hu�n3�a���a�+%fmߢ���μf�DZ�-����]��M�Z�T	����l@�D�g���{m%%D*B�۰�i2;GC߂ڵt�)
���P���ɸR;j�-8BL�1`㛺�9�Z�N�#���J�Q��t�LMw���Â��ԑn���!�Hȋu1s}��LN��^X�bn�� �4���ئ��u�q@a=�mu0_Y�( �DF���.�e�ewΰ��|�S�{2�O-)��ؿ���|��z��_�y���v�
ŵ�����l�t�f�����~�xv�ڊ|3�6��Y,������� F&�Y:ٗ}1kʞ
,{�2����3X9�۰=�7��p@-�S���J
i���+��j 7�3M�������aC m�]<����S(��+1��.����ޚK)��*��H�U3j�R��ށ���s�x��|s�ϟ�3��ʤ�ƞ%�5��D �� ���g��n쐄��Q�v�n�3[��Y��!����ns�� �o3��֓@|�(��\Rc�!+�s�[�!k[�r@�$��EFB��@O�T#o7�lJ���MK��g�)N����tH���[�WmP0i�D<�6z$�s����_/;!6@"ߕ��b�<��r+KW�l
�ޗ����	'6��3Ǆ^+����)��܋�����	�ԗ�<Q���.��n�;i.��d���-�H���!^��h���6kDRx���:<;���$� P*@�����YJ�y��ú�3:Q��ĭ]/������^4�K�#\N��-5u	�h�*���R�# w-%�)��گ�߫p��͋�[�}�H��uf�i�8w0A�m��y��]���{z��knY6n�1��7�� e�5��l ]�a��7���� �m��)i���]���b
��0v!� , ��sXe`���{-kI�h]�������O����s�=���ե����߆���\a*��1*�Od�����{�����Ը��'`B����U�h����Md*ҼC���C}=�~��������Z�śQ������l�H��-�1�M�L�5�\��w��t�Ⴔj�5���T,ȭ�d(�>�1�G����� ��nR,�bS�:R��F<��.��7o�$��O�_A������ � ;)F!���n�B�D�F\e����VL��r�gG�C�S������)g���8�2Zvؚ$n��?NG�������"��!'7A�ZfJ�Xua>���-���`M:!ck�U{��!�/:��q�&sc�����B��������&g���օ>��xi�_萆'����m.��Q7�}�)�QL��؛ӱA|A����IeHN���o���e��V�z_[P�-����:���Т'W�n�p�����Or�C�m��.����}���0�g��!���^��i��8d"�'�Wj�GO�����,4>$��F���B���4��֫��]C��i�����|:[E(:3�c��8�S�#�/V�˟�OYu�cc�=KA�R�0���b��)����^WR�D�e�$�Ȼ�c�*b7�c����Ȏ�]�Yګ�r�9��������^v��EG��n���{��J��D�,�
M	ao`2�8�=���;7	r�H_l��T>�+_2Sq��>d����,.2Y��Lۗ���dZ�m�SC��u��r����w����^I-�/�^�D���b�<{+����`��\|��D�V�'k�c���T>o������I7���Ȯ3T��u�v��x3�h��#�?�R+TZ�:nD�9�D��o^����1�c	&��Ĝ��Hq�;Io�A=`��T�&"@�|_y�A���Co<������~��
���܄1���Š�D��y�+ߊU�^�s�o@?���G"�;���9�oH��8��$|î�=��ǌ�f�s��d,+
�ܜo���<���F\��$�;Z�� ��wq�-~8?� 9c�݂����<��xB��.�� X*N�B��}�����z4FR�?CL�B-��g�7�Χ�1�����sE YZ�����IȝG�;q�Dm�`ظ��L��U���w�N�J]���@�|���J��
פ�~�Pp��۟����_����2$^���!c�M����@�`t�'�q^�sm�`�&כ?dno��4�V���]������n�1p<��m��� ���c��0+J���������n�zڡ͋��>�9�M����{�g�wIHzK@�9 �q盖�I]1�1�oy�N�e9s�=>#�Z�?�l�J5w[*D�q�����;*��-��7<��;����M~J3[N(��b�Z�ο����Nm>En�Ru�4��sy����`<��` �z��m!�����ﮙt؊�H�r;���M͈|�*5� I�]������k�+YTn�VF:�4'Vl�T�4s��/�ec�v�x��M��'A2���-�;{G�;{�w�<�w�-&꜓+9�b�1���p�A�p��7EV�z��▣�(O����*lwΫtK}Ô�����~w�"k�Az�z���ݣ��E/vE���v0�����؋�#�vVб�W~�rF����C�I�_���:y���h>N�E��DrO_��J�5�A$�rlh�%OO��-��f�����n	��&oJT��:In��f{�$t�o�k%�1��NšNMNKՇ��5���Di�=�)�C��iZ~���c���i��K�\�dV����gK���R:��l=f+{Iwy��'~3$���? ��ML�[p�yO������S+��l�4k��v�+��-`ǀ�݁�*�~�T�R�yR����eE���Zv�Q�a�V�y_��90�zLvM�Lg������]��a��Ų��b>�N��c��PB�!�,#i��{����bÊ�;���S��l�dU�D{�����f�.�f~�?T	9vJ,yP`��t��7p(H,��p�?{�6�~(Mn�~]hQN�+2�f4S+�+�3.�N&����ډ�z
�/1ނ�U^��N�l��v�`��^�,�8����f�&����#�5^�o�e�P�&Pz�Đ쇓�%�D;ڲf�/��mq��D|��j'x9��{Y���m80#�	q�kF1����e�NՂ��>�x�[%����� u�1�m�	�{��$�걏ݡ{�5�z֥�	��,
֡���T��f7��a` ��e�N)C����vQ��EN>���4|��:�2Ө��,Zu���ZR����u���)p)C�1!͔�=�~)\�-`c��H�,+�r�.#6Md��������o����7��l1�����d�c!uq�Tnk\el5���[�>f�P>���(V(�ˆ�C�EN3�\l���yD�e�f�s-2Ȫ���]��Xz���#dp��	Fѫd��u)�T����O�Z%)�݇H�`���I�C��_���$��> BH�h��'ur�Or|[	���Pk�������S��va�/} �a<��*_��?�!� �ix82s� ���v�7E�nmz�3�)4.����^�����\� =К�ƿ�V��Z�.����!VY�w��c{�^Gp������Z#)��p���䙹�%��o����Ϝms��q�Z�T��hQ��r���R���c�j���������`l�A��*��::��ߣ��g��+y�s�Lʌ>���!����槻�O���.��v�bY��4��
ڮ��k$�k]�4K���h�*�Z�u�<��h;��k%ө���<`[8V��+�qT�_��}�qn�fGGaf:�U�<F��Nw�&XEs�;�/a
?	����L����8a��q
�ت��ciJN�����a� P�M:e��r<�����w�)~2݈J�~:
n[�	���s�����)��֖�R����bV$d��'��&K�]�l��SP����	�����y0��o�j_yi����q��6�n6��:J�K���p�XI:���zr�v��Es�!��O5>����������Y�>@循��Ǥ���}�������(�������Sc��K�_$�dH�[�|wt�Rl��"�+*��^��Bi��xC�(Ņ�����j�)���"�����z����R�f̬�H�l�m�h�2L��Q>���,:���LF}��K_ �)m��?`X�,)����C~�גO�'޹�{�U<=d��D�=�*��{݂ԁH�v��"�BT=�5��2<Lāj�z�{p���Z`��:���2�h�%���z:/걏�L!���/[j�y��t��?"���r�if��\8�gݽ�F����+#���>�2g��Xf����~�� "�9FWئ�[n�� ��2�kZ������,�I}���n�d�`P�y P h�ؼ�p��$}'�Ҋ�ΨbS	=�N�9��o������I�#�&f�d�N�S慇e���U��:X���#�o�+�K(�f^��RK �M��t����p=��.}�b���`��M	�NW*"�����:)?q����g�=�ë=�4w�9��QaN@��z4��]U�m,G��5h�ěxu2�C�Cxd}��8�c�6��C��+�V� ���Q�˽�b�y�0�3�	X8��(��<�X�<��L�z��Nx��[�x�mw�7���J��WcL�l���n���%f�[R�
��.8��x����9M�
)~-Z���13&�t{�b�I���q���{v���Σ+i]z���y1�m�6�'�!��k1�'���%�r,�#)�!���:����?���<ޯ�,K�;�U�?���x|��:�ܤ���-�4@!_�+0���ݺ w5�v!���s
,!�E�VB�c��dse�q j�<��ͱ;��M���\9�$-�a�3@���^-��B����2n2����u����9���4i�d�&4Ee*���!�!�U>�_�F(sv
פ�0�['q!�8G�!g�v���
�� �	l� J��=��d0�'��m'b#hv�		ρ���e� t�������AU�j����Ց�vP���I􈴁'Z��K�����_� _��v6���Ո�5m?z��
g������!o���N~��hle9�ԡ�~�������Cy<��0��v���[�o�&���4ܰrH�é�q"J�Ӓ3x��DF�X��v)c6�>�kF��rr������ ݻl���9��һ1++��L\�ž�d�G��q6��>;����3A
�3&���$��M������2�������T^W���f};�L����y%p��盪`!C	Di%����H�F�D��d�^Z����Xyk�$����䭝� �k�/�2)�`�.��	֑���i��+I�xo��m�6N��_>��+~$��4��r�d��?��ڄz��rZW�ɜ���I�x���y�Q�̈&�c�Q��@!$�Gm����Gz?C{U%O�N��)��B�����	V8���1H������#�yK�����.�#��}��v\��}Ny��7�0l�����*@��r5M��hH�0lB��R�� =�h6>�^���y/2��ΐT@[/����0��]��#�cc���	]�r�܏i�,�LnAE�**^$�^��<9����3w'�GT�^h@<��B9���50�s�
Ç����x��ٺRZ)�E��E#o����K�=o��FY�W�T�
,�Y��l�ξ[n�°��05��Uy}+�6�"{8��c�=�ڶ�i�}�o=��{� �E^m�B�V��4�`I�����ꮮS�wl����]k�'��[�[tSzH��^�e{�� �Z�vy�n�Dl"g
�#ަ	�v�I,˅Z���|\�ڙ����w�uv f�/#��!��G��U�|p�q��Y���[Ȑ���8�Á}��
m�]��ŵB�P@XY�Z��%��w�4�(�p����$l��e�5Z���q��lq+k^]���u>F��٣	5o�'�4����t�S��C��.2�NJM�V��%���V���Eo+(�V���-��5yRn¿Z������H45t,�V'�9>=�`w��kjobq�U�������VֿOA1�2�6v��?`l�+��p���0c������\��fuw��X�U(AT����O��Di�g�r�rjyv�
V_�*�7�p����+`�%���K���8̗R�'Ғ���pM�ލ��K)M���x@d5�˨k,�_E�GdiT��BA�{� Ͱ��8�������<���ׂ���rf�g�_C�3{*���^��TD���LEɽ0�'�v0FIS'ϫZ��'�3?�����%h"���������R�����J��yk2�5NR�� B�8�<��wAKY����3ua��Oe��R%��3,�sq|�d�h�љF��F���z5-�&����G�ED!p�K�`F5�s һ��ݮ�w�ϼ�X�+a?]����u��u�"j��Q]�)�+���E�?�b�0jd��fZ�&[hC&��O�/6G�#D_��� �����}mT`�9�:�,+�7�I�I�&�ֳ��|�GA�_����m�5(TE�?�?94C���y�i�$BX���^��1����Od�p��~�(��Bֿ�,�q��4�{�w]���N�NxNN�u�;��P���=���_�^&��w�,kٟ�;W1#��M�΁ק*1]����w����.+��+u��q7/n�Na&1x�.�x!*|�mI�T�����a*o����.��8���
� �:�c������uT�G�s�e��T� {�?���k�e��osAbΤi�bL��p��j���=e��~Ƿds�E�X�������Z�m�*�Z-U��)j�|x+YjMCU�U�@��6�x����I)a.�l���0$�T"=t=�D�������m%�<A�bi����[��ɡAp^¦�����4">��ʦ>�ڇ���ǐ�DL:e��-4'0�
�5K�ը�'������pK</����I��1v7|K��ڢ��Q�sI����x�	iP_�%��ȭ������� �Q��_�?�k��"(T,����}�eK~g�	2�D�ï��ǩ����;�Z���������:9uw���h�����UR�M�Bhp�m���Sb�B%Rlp����J�=�W��n3{�8��-&p%�ϻ��֡�����Icm殪�lW%��@^�6��A��ű&*��'�w�94��wkL�~���±�\-�P��&�(�P�֘W��;�W_f>Bw�:0Ŭ�!<��L��lb!8��l��j����X;ߛ򺑻���� �Y���W&�k��ĝ����Ŷ�N'G';��q*�_Mi�bUwB�K�U�4dE�:W�gd��|Ի�G�sAí"\������[��SX	���"��%�G��J��q���!"w�V6��vNߕ���̹<% >t�B��$�)�\�0�W�4ґ*%Ŭ!݂�F(�Ԟ-�/��2�!�\,;P��LE��ǻ�1��3�X�q�Om�.�En�t�$�g�.}!�Øa��&��X�1�����<�mlP!؁+��)&��9q��k����V�P:Mw��,��y���o6&�l7��]����р���y�f��Ϯ��r<~A�$�������(`@�E
؅?̢pȶ���c���E��\!"��w�^>��)��?��n5�w���J��jP�߾����o�BT�Oe�@`��7/��	��g�Wi�1���|��ZЛK���4=�'�W,��}��e2z����Nt��]��+��n��#� �	�=�ס*U�{��R��娺:
�D����m�*��?Or�l��0_u���$��'ZQf�lG,7� ��XW2�����/�8�0IlTSӼ�F_|<W��
�}/_Z�<i"&����&tu�VÊ�FDbr:�[�o���[����l�\H
+gz1��=A��L�'�mWN���d��л��P]�r�g������Q�(�h�"��f,�n�"/y���J5����[Z� W���ޥ���NF�'�Tq�5�a����ǩ�a�]Β���C�.{�COn��H7�b���P	e2˥��8��W*�d�%���+˼\�3a��^��M�>$�(�(ꚁ��r��$��L��f$���t�����ݯ�<%l��v˞mK����K��m��Z=��]pj�
!�wc�9�("H��`����lV�yŝ���؊.��RR&F�C6�kO��a���c����a*���`c���ٮ|���hǈ��8�p�Cs&aA�O�.��PD��`�B���4�$�� �t����l�o�&�|�ߘ�(�we�08@|�7.�h�X
���`��o�i��\"=�{�W粠��ޙ��	W`Tf��F�M����Ko���������T��us՗qu�s?��W��Jz/h�������_�x:1�#u��� LL/�ݱ�#�T��a�@WhU[�C?x>�O�P@3�C[h�������kb��h��~�l�d���0\MpM@g�c{�P�K��h!��6�,\-��d���	��V>�6��
��o���9��ُ�.7o�1��ͣJ����/���G|0=a��.��ɸ��	h��G�?Ty��y�R!a:B[�P��l�˛Е��F��k��oX�[��f�|e��m  B����t�CmJ%� /aS�E�Z���Uk #����ኊ���Αi��S�������
�|�	a�3:G�T��)=�X{��u�2.#ɉjb��Zy=�$�e�SI��@N��E�E��ᵺ?�%���2	���#wK��A��$��ڬ�]�"˛ ��LﶾL���KO�)��'~G�������ɪ�� �>oVEqt =Ib�;�q��!^�b�HܚT�0$p|W�	C�&�'L!�:����;3�Q�iӔDa��?��l��j����;�е	�B2-�-�Iaφ�vN[7��}-s�i��Pڕ*����2@�':�"�E��c5�J����ϛ�d�'���q�a64�Jio�s"zY�$�Q�� � �ڽ�]�
4aUA	���&Vn��K�����Px�~��Z�P�T4 S��`3�+��n3���}�c���{��m��.%Ў{����}]�ȱ��bS�pɫk֏^B�:%�}�'�ř�/���L�m�ͮ�/�pGُ��P̖����ʿ�3��g�k��G&4��aWIǜN�6$�߅��{�Q@%h��#C
eE|�ksV�`jߢ�d�Sf?�urT�ԑ�!Q�w����i5OF"��W��I���B�V��`�`l��T���s����2,)�8�ؼ���bY�jo$��v��V��&n1(ⵤx%˷���/�C�d�_i�}ic��^�[��{;���}h7'�
i�Gő��6�X��ac5Q����Fp�#�{�%�6Ew����*��
��|d�^Ԣ���i���k�m���A��̑n�K�Z���9���p���շ�5��o �u_�8�r��t\�hI	��F+���D���eħ̡9��e6㱻[�H\z�3��U�e��Ƴ��X>��{l��-�5��eܶ4��^�ۦ�byV7FY��3>�n,la��;�Ȧݽ6�g­}��#(j��d��ЛO�?c>���OG�Csa����ns{C0�זS�w"Tt���W�;�dHI�2C�Ut,4��4m1���f�����	�v������a�$��;�Xm�� ���7+z�������g����[��#�q���$�:����4����_溻+��V]u�M�$�%����fm���BQ4��X�!ާ}�R}�완y�X���^������o�@\���d`G�z���{�{��d�����}?��J@�j�+we��)��(e�%�Po�e��>h�E��9��P�T�~hS	*!ǵE���u� x�)��ժ�8~�qv�b�t��A� U`t����Z����5+d�u��Ò���d�ٽ"���Ƨ��Gx"���B�4��0�2S�I"�B�1�2�穕(ua������B�N�Kգ�xu�=�8��rs�@�\��_~���[�x�������g�$kH��Ă�qؐ�!N�B�f���jz�#[ ������w�T�������**
����1�W�v@�{��Y/S�Be�ؙv���V�f2���ʅ��=0㌳���u�u��x��{e�=8���Q�d�V>���R/[a�Pur�m�v�H�w���n֦�/7nf,B�`�@��u����s
�i\�okݟ'D�>��aD��7�M��_(�z��K'�v�I 2���1?L�`u6�͗=Qā���|E�F��)Z��f�E� � w8d��~lII��f���YsI�`#ac��T�J�@�$�$��F�Y��u���-�|>Pu��
�*!���t�( �:x%M����=G�;3-���+�*�_�\�v�V�m�?2�[�Kx �7s�l�]�!�:~B�U����#��rc����� -e��k� 	�y
� 3�]��b܅9hކ��{nd��y��|��gB1r�qƙNn�H��C�pgS+3D�뭯�>tcj{ߺ~�o.x\68�{��i ��b9�tBoO�6P6�fɋ���Y���<FH�?D��#�c�ߑ�� = �_�U�f@;iV�N?"v�RiTr+�co�Q�E�`ׂMk�T��*�:�@�4��@\!�N$�U~�?��[���-H����&?>���\� �p�fA���e�m�	 -��r�±�'��UA=/���|�2*�bM��9RJ 1=���~j�ʅ�����`)J	̳�XRVH3�u���48�b9y�̨�pҚ�1�!���e"Қ8 䞄m���_aX� w�#{jֺ
F:]&��*q�&?�|�X|�T�(l����pon�^]�%a`����1�;�K Z��ڕ�:����zU����r`�f��<�����&��{�s[��k0���H�-s�:��4�5Q��M�Fţ�ɫ��-w5������w1��k\/���8?f-���QV��#!��u���{�d����K���+?W�Vb4�Nɥ+w��ر$^��e��|�[Yh�ׁ��wEgz��`\jM���8�<��L��t�ڪI��6�S�X�N��q��U:�ee�cWV�y�
6v����l��Ӹ��[�9�g�k�+��J���g4���=8Ce���IkUX�݁� �
��?%5P	�+#8�̈́�S��(@.�^�*��<�X�����#���J�FJ��	�C#�&I�crMem��Ď����]����m#1}S��J 7����P�a��!�5���� x!�YU:���"+�`z�
� mh ,&|��q���� J��X�FH%1|�?�F��0xn�
�W/ܳGT-��,C��ӳ�-j�7�af�
�jL����[� ��Q>+��Q9R3J�����H�u�7�J�j�/|���9U���ӓr$�����Пܞ���ݥf_�A�E���EF���\_{�'6/1Np���]�u+n8���I�t����;6���N�%:)�8AE�j������!��G�0is���lvr2��$����V������Q�~'Q�C��9O4iMԎ��J��6a�Έ�����Aqs�}k�_�V��(�1*�D��� S(2�f�Ȉ�#�-*6�M���� �Áy��I�s�-@�N����-:��0��� (u��H��� K>�X'bVY���U93���I����ξT-�����Ɖ�V:KP���by�.K��r�Ry�ʜ(�b�m��r���A���+,��'�qRQRr6��@K����	�&S��Fm��)�L�Z���V�8(���j�1C��/�!�����͵^�t4�o���y�I~�%k+���l���A,�/NU Ħ苖	���[y�jN?���h�u��Cx�B6�'�Q�֔x�4ށ����2S�В�#��>�?�U0�zÍ���ÙT֪k܈ه�����B���<��1骾�܎�׿(��L�W9��, �E��,��#`Oőv+��X$FL��[ۋM�S�Ec�!�*R��[
@�=��s珖�����Dm2��~��ɉ�1�n�^�};��3�����X�Փ�*vS��/N�0��̷�z6����x�clØ���0��
Y��_^]��_� ���U[�3��^�,�,�?�"X ��!��ї�c�f&��{��oFg�փ}���n���h_��)�"�͐�o:5��ѱ
��L���-�$۳��ج��<�.���Z�p��2�2w����rHz����Nkm�V�*�F���.����� ^��b�Vj5��P;�����K�~rX�)/b
)�N����X5/��{	�O���UbT�Y�{��L,7$ds��1^�|�i�T�61���B��>2ӭ�� h�V��lK���ո��wS�Dtn�x�D�w��5I dDK�c�K��w`�2���$�}y'��mr,��2K2��=z�|5r+[���Ĕ��O�夝����Y���(uv�a�*5s`��p���	_��S$��>9��uQ���/5���L�\j��_�v�R4�2���7oz[�TA������kb04��Q����:m2�3�^ܤ��w2��8�Cy{Q%J�.��!���ֈ�ۼ5���/1�&�3��:���׹�))�z���Q�~��jΙ��6�t�0`��ĺ����R�'>SPM�#��rj��k-QVZŔxa;�#I�
�� )azy��_�@͌K0�+B�H0m���W��0��_�Kk����RU* ��J4"��è`����DN���O��������*w5}�Ԁ��1��Ny	�ih#�va�^�R������n�����1��P�a�ߙ���i��z�r""]G�NI&��YS�q�5�2uY��ޝp> �XT�n�Xߺ����\���}��uҿ#7i�w�J�1�:�<De��>Wc�n��o�����!f����B����c(���d�g`o�|�Rm	͟j���ʹ8�?��}S��É�7{۵Uv2�7�i�Na^�[:��/tK|ٙ5�M{K�x{%�pyh1�΢I'���g)PF����@��Ov;Wx���2�s�8-���#�����p�DX��)�o��?G���c/���۬`c�Ǽ�m��>笹Yþ#mY4������?.y���(��X@.T��|��A�,��V¬�b����~�t���F�Bp�g,GH��(Y6nJ⺘����?#�?��K��-��E�E�!�ia�)1f��&��٦R����X�h�]�pT�p���*�$��XQ-�٭���i�G�����)�"֢[N|-�;�	�.*i32�h�H"B�����y�����ED3��#�ā�y	����r������]�Dv�M���6O�|�� �i�4�;1z���+�G�D�K��:C�ݰ��8~10�!J����X��L��� <�/���t�(z�A���9"�F^�키�S�$.+1��ٙ��DJ��B���f*l��q�[�8�v8.�G<�i����o��58��6�T�t�D��QϬ�MӛB��sx��A�4u����V�#`�|kmJ��u��:�q�lp;��?�%yv<B�L3�z����(�C�T|A���'+�V1!ߛ��t��-I��P�8<tG��d�0���Y��DݹT(� ����:zn\�=��F��M��$�$�}��񬴭�To6�p������H�FTL�\_u �����2{�t3�ã�^:P���`Xv�7	F����^)�7��3B-m~�]Q��Ap����'���4��8�i�Ͼ�RVח"���D_ʰ��H���u}A��,B����q�9�W롽�.t�st�z��0ꟲ��d�[ݏ��wQ?>�U�`�R��&�'j��.l7ϣ���t@@�Ј�7�%0�yW�m�i�pX��J����[p��{����#L�NF;#0�{2�e!Z�J? v��z.	�d��;ް��<TcV���`�P����\p���}����}>��ޜ�y�9e�qOR�ǫt����aE�՘z(�%�[�5�0�+��E����ǟI�P �&w�1D!J�VV������PDʶ�*���J��:������E6,l.>QJu�V�E�N��;�jm���b�������㲞�*�n:F�쌋�r�v����cdB��c0��������Z�9d���!�@pwqا]w@������6��5��� r�a)�3�b��E=���=5�je��V�)��Kt�G5&Ls�>�TZk[ܬ���;h[����B̎:���j�� +��	�#�[I�Ǐ�V]gu@���m̈���I6*���������o��ad>�|f
��Lg��\��#*��3]ϧjݞ�¢@f6��+O�!�J8����AQz'�8I�ms��;���s�`_x��m��Y��C���nm�;�ܸ�9���{���|�]�oC=W��~lU)�8��H�Sٍ.�[����E��J��[��)!�:֚��a^YO	�����U݅>gɪL	@��ۃ�0������ˢ�R��̗�����(���]����]�TdK״4�9G̐x�1�IV@X��Y�������~Yd��%�=��P����9�.��@�}	M�8����dz����T���a��fk�;���6|�[.縕.�·N�t#��П�_3DOT3�	��k1Hp+����f�	�-*g�����\���_�x?Hr���
m?�id�GRw��W۷�K��`L ]��J����)R�����ԯf��i�ĥ��CԪ�?�5�M�^Vq&� ����9Z�Y���mR�I�d^Qnڵ�b�ts8� |U�ɢSOv�Q��v �o٩~vά��a��YV�d
��6�3^��+�94�ڀ�D�q/�?Jb5ۊB'�e�?\�݃�R����`�f�a:o\{�R�_�}Kk�\��s�MAޓ/���L�n�3��^ҍ���8Z��a%\`�u�X!a�kzQ�l��$�q�u
n.��.Z��R��IfhS�GL�����f%�1d��L+˹�qi��lD*u>��1�ػ`�ߛ���(�شN�Q�7�bN8�V�4���9ns��W�1Z����<A���Pp��y��dEx�N��!���P�-�*�����ĭ�{�����NOe��DU�pP�3+���Y���p�W|l'�_�s�[�oK3�Z(���w*��`O"�����EzwSBܩS�
�
����J7�]ڜE����T���`2"�Z���0)d���n-���zM�`z>%H���`j�loN��⯌Ļ(}�"�pk^��k���
��}�O�y��D��U9ݘ�08�Û��{��L=	޹�#k�4e+�g�@�!~��?b�rT�M���=_���"�P���[�<�s��VN��aж���\�]��гx��p�u�Oxv�Iz��6�ˎ�iն/����Jt�t6��v�#��u/v#9�Ec�^���,h�������8(sWp��)�4��C��A��Q����[�k,4��$����w�������βy�0U4��_�'��~#G�����su7[��Vn��傿0���t��b��2$2��zWF�X�;���E�a�_��ֵ��0 �T1QT�W�������o��f���_���
F���i9�C-�]PMLy�W� +��ա��N!�
���jQ�˳�%� 29|�El���.��ջ"�^���%6��5�w�D��2�\�t�j;xI)�/\U�M��+J3Wg�<�e��k�a���ץ.���~��K�\_kJ� ���td�bH�iO)�8���ܖyQ��d�g�㷍��(��*Ɏ�(��=N�����fЃ�F���X*�]g�c�Y�)*C7����b����� �-7�F⡅���  }��c��g���q�����b�i`!������Ė$�%R��4����R#~-�? 2{��^ �Q�}9�Fr/܀��a�!����L�q�G��4ȕ���:1���.��
��^cp���ZǗٰf����^�>�4�x�B�U�GQd��(`~���JF���5O�o!��j��U������0W&X�g�h���pSƂ"�M7nE��f�����H�2���y��Юp����6�
��)x�ˆ�-˅����.T��l*�1�,$�P�ѻ����&vj#y=���U8(���� ��U-�������_��28ŷ�9��	lFKڀ��J����їʎ�׭d_���t�*ia��Xڱ���<ў�빼m��H.a�P��oqg�~5p�/o����W��qYjIH����N�~��e�Y	�������g:d�2Z��L���~_\=#F'Ft��`p�U��Y��@�.��7�Ls<C]��M|	0J�|ʽ���Y�[�J���:��3�"Õl,�qP�d)��d�����ǐ�%Œ/�P�ӕ�[�Qh�8\��m�k�ש^�4��a]��'bo��|��ˈs.(��+�sF�K�X��i�������Z�d�N�n�-�,������)?y����P+�O��)�Q��bhM�2{��6F.�ur��e��9?X�g	��;CX�qE�$��Qě^9���s��5���g�8�ah�[9�`_Lw��8�O�k�^V{��Gt���6��P~_�6t�򭆌����8*�zaJj��W}L�� ?;>��o7��,���0շ��	Ɛ!�Kt����]в\o=L#]��㌯o��\�Ha�C�!���LY���X�x�v�Q�4Qs����7��1�_�^��ZM�y)h���vD�,O�i��M.U�r.]d�*�>u�'ef�ED���gf�8je�-�6�R[�?�u����^}
�[YB�m�t?�:�Czs�����)�h����@d��i&Χ&��*9|��o�X5�/'6��Cv��D��]!����� ���t/r)����IW�[W4jU�a��ˎ[�h6ٶ�fᓲ��_��T)p-C<D,�=�9F�UaV*]Ɂ���q�3���7 
���讀\�)�𖏟p4Y��*¤�3��Pύ�L��▜�~�R0���1j��%�I�ä�6CY�ѨM�}t��'�0E��*|GM�v�����b��7���cM�|��x`F{�M�hDv�S��ȸ�����;��}Jgmҷ���'�ҁxku@��#�s�yH�� A��Y�a�4j���Y4��Xg���A�,��@��������g0������)����;C
�L��8�h��0?8�Rxv�yNh�:hn ���-�pT��Ի{�M��Ig���!͡�&�U����R�.�R�Q����?���WW<6n��J�^'zNv@qk���JZ�{UE�ʸ����>>;�����f����ѧ��+��T�QO�;�Lo�D�^�l?=0�)���=dN��|��}C0��n���/��t�<WF�G�,}#����M�wʦ�4�'-lt�A�����)+$�TEFg�m�$���m�|�Jh���>׏dXv%�.5�&�2���\tT"dXR*e��E��!�@�bD��������2�R�P���ÍT������xО���\�xϙ*ѳ{�8U����\%�ɮ��.�v�K^��9��M1ח|f��j�K1�TlB�@�"�z�Ʋþ���p)ۜ�wA���i4Y�60j���{Ó����	�G��H�B-tS���/0��K8pTշ����z�����c���i�DP��k7Bȇްw��;�%�y�"ے���u����_��TQ�:lZ}��E�d���7UF@?�w{����Z�n�x�Z�xN��JW�����$\ݓZe�I:ɘ䇁��/�8Mr~�+�Pl�WM� J���S����e�[�@�����8(�T#ƽI~h�l����R�3�*����#b�L�
�6a k�1X�rP9h���)�1������7�ޝ�O�l�~D���uZ$3��ˀV�h�,�����9"慎9D�F$�d���E9�U����9�gY�\��✄�n���6��8�Uf?�Ѭ^H��!�	g,�Z�Wݐ��j�͹3�|���|lC���8T�|>��A�>4�Y ��󆝕�?�^թ���x�m�X���2��s=Z�Z�<���4�����xCx q}Hh�J�Q�`"���iM=�H�n�s�H]w��6/��)^�س�u����W^j�+�v�N��srƞN�'���{Ŝ�`���!P}���Ɉ����,��OfI���ʍ���� �8�ضj�F��1���5����sVS��	Y�� ��"��$���N�[�V��oR,ɅW2J 
��ǖίeN�zĞ���dz��Y�ɤt}}x;�� �_t	�X��(	�c~JҐW�$䟙#�k.�|M�)��w��M����W򁜿H�d��KT7?N���W�T�;���x����>���&V�؂�c��<�1���P��͌�'S�v�)zB��z5Fk,ki���;E�n�=z��*��d��7���a���$M�@T�> �B���z��v]
�M��Q'��i\���9rZoƷ3�Q������P��TIi�Y�4�)#���e�����;C5�~9mu�� �n�v�*9���X�g׌x���_K���PuY�,��}�"�������a0�����yi�`H-+�г�U]�o����Yx_u��M=sKH���Rd4�>�ɐ�ӥ�]Q?rs̓Ԕ�i<#�Rs��inyP���`��Q�EGh��ml��Q�u!���J�v�?�u�'0Z����ԇ�4 ���Ǧs�9']�]	��SJ�F�b,��XS��dc}K�9�h���Q����8�F��0�*tnSu�-fp���R�������ٶ�`��Em��Q�*��
��N�-h}?�p�$�`�#6�w������9��&ߠ	�k��	�?(�̈́N��L�'��dH5���f��.�J�TAT�h�W�_�?=���?qb�x*'�0<@��6�б��Η��1+ʫR_�*A�퍱Q����aR��!z��p�/	A��i���W���#`�-$U�����wB�yHkNE�@��PW,���̃;����73 [>�5!�]���d�og��ë
n���,1������ܬgN�n��Y�Fp�%(�Y�����Ir��+��!T��30�{}F��+���R�ԗW�q3�;-�M56'D`R���hL'���!|��7���T+�����?����VWyf������4o�\QI��J��sxj��s_ޅ?K8��n��ҍt �ORd��9E5*�	���\,��b�x!d���ю����E##A�D#��(�'{��}yq�M)-�)��N���l"@?b�-V�W/�T7���ɇ���\���r"�� d��&�b�b���j�͓���HI쩫pf�YVr+���H7#�����W�b��>����3�qX����
ԏX�D�c(H�~�nR�E��~Q�!R��1!�Ĭ
�d�'7c�8����S�A���y]�?¦㩰 I��O.xKCE�H��=��>�R�d���ވ��� Ie��!vB���ў�Z@)��B�o���J������3��x�Zl?2=O���+��Y�q�ȴ4�|�i�k�u���u��F�E&(��98�D~�#��ޒab�bS�������"�cnyu:�[��&������$<;��t��.�"XYd&� ؽ��nH$l�cJ�����>���"s��6W��8�����RD�t�3��?�d71D�R��wp�c��zxW�yO�Z�Up�Ɦ��G�̉�;3	?��5��Y�CL]���xL��k���S�T���x��ṭ�NX`��Kp�.��%�h��K���!$ʅ��v����UP&h�¤�Ѝ:��􉡶;d����������M�<��O����v�(�tPv���	�L�Z�J�ܙ�������,[��:����:�Ì8�	d�}Y���|h~��	x��h��^l���5��/��*N��޼�CeK\�.�ab�<o¹ �2�?�-�ڌ��4,sw>tk�`�(]��*�OYG�ӥO?�A��$tӖr-)�ch�̽J���]�����-�%�8�t'n�ܞoR��&�ҕ�ǃ���햨�}��<i`4C�e��'*�[q<HH~>WZl��`����[�]绩<�Ƞ��% �hWv��C&w��y,���!�X�X�P�x�`}�?�)�X��.f�c�8ɟ�-`��^-����;�1�Ӣ|���bB� <�Y7��V-9�}�>X���W˯ .��}������A�mg��*���O	"1C�!2�f\��2
�5f���#�&v>��'P��IC��Ba` ��8�mI͖ �j������I�g��I �Ɔ"M&��t��kG�����Ͷ��Kz	��":���DÄ�"VX3g��烠/Yj0G��_�3�f�E�g���}A+LB�3LeFw�<�	X��6���˝��]Z}�v���'��m�Bb����'C���}3򵇷�|Џ��{q|�W�B˲c^����l�!���.!(����:SkNQ������)aA!�]�?u�+w�-,Bǔ�<�6u�|�@K��rn�25�U�\�&�Q/���/c���5V�_<x��g�)e��M��/pq��������i�7�ݞ�ܰ�EM+8����7�1,[�L_&qD���,�v����a��[_��u޿)4���,Ǡ�g�d�IF���W�q����_$v�q!�����qE����A��q�T�����~�F�Z��3���S��
^�0	&�#�y�0��2��f(_�V���<�'�f����W#9�����>i�X��<���r�K�}f,4ri�na�-���:��^�J�.��IJd�"�z��)D��PQ��äQsV�Wt�e�+ɮS�?�ߥ��cP]ܓ�ЬO����RY�M��}��*:gT���n�qsȾ�l���w=�$�ϕ�}��U��. �DY������uq�%uc�J�����рK=} ���_Atq3`')yȜ+TN�@ϗp>f��e8�&����'�lc	���f����>��z�ls;�|����E�G��ǆ�l���_�:��'g�v���gt=������bI,9��`RE��W�u,�w	nxz�惘H�!l�*��f)�}��^��q��a�]���Z��[���;���W��馗#�دg�f�oj��_�~CѾ&�'a���t�A�Px��K�����M����W��8�`�Y_+ْ���ź�H�#E�4��"�4Мsl��i�~|�5\Ch>���$��-��%�=�C�<1���~`�9Eq|�@�d��!�1��;OR욚'l�8rop�-�i��#��y�ȸS�g�C=3/RE�0D�:�>��w�~%���\lzYw��a��U����R<㳻��#k�;j���\�/���2vE�����ӣڷ[T�"�7|{0�5)V�2��7��"✊Twp�>��%�W�� ��U�������:�9A(������=M����Gs(���9��Є�J�v��U���01N�A���ǹ���{���L�q���}�������i�X,.ZY]�ʶ����)��f��qX��+�հ���&��B����b�,�,r���6%���FI�'��/H�����-T�R��
p��a��A�D���b��Y�������~H�ӡd���=Hh�+�"Ef3U�k�t�[�0��2b��]/f�.�dL5{����5H]T���n�������p�n���e�S�潛��4�;�pO;^���n��6��K;�KVV�JP�4���[��'�F�$G�t5%����Pkk�êwQ��>�$s�c�8�R����W���[�bݲ��'S;A���;!��z���nj����N#�˶q�7�W|�ě|���.[*7�����<F����52�]�
`�U*6�ؐ{�<�4B�卌�k`������HN3�T&�Z��B�p%k�߾�,�ƍ�u�J��Ac��F�?��>@=�&�-�@րhƨM��Y�҈־��U��ᝤJ������j���%m�c���UsH��ɺh��Gul:Έq�2
?�+��mvh2� ��2 gX��qRY�
E�g`�N���7���e��ڣ�7��3�`�����q`� Ȣ�ҺO��g5G�Ǻ��e*��T���Az��)�:>H^1a��ڙ���\�8����9�	�Pc�G#�Ѫ�^E���>�𒽃B�m��QF ����m��D%�&�Y�n&㠴B���#�
����Ԉ�Uc1�]��%?�s�@�ͪ��2�:�Z���|U����+�ᴤ�7�a�e���Px��<��٤C��Z���Zi�j�zx�P��}�j�&���.�'=�i>>Q��'p`>��'�����`Zs�(�%B? �>H�5թ�'�g��;^����N�nH,f�.��+!1�<�JlCA�(�2�;�_d���}py��4�eG�6/�S"�f8H<�r�uyT�	�(p?@:���)hܶo� [�ae"~6�i��8�c��o'�)8����B�8���J�1���Ϯ�K���">1ke�^�3�h�`�������HO�W�������ؘ����ఀ� p+�������@-@��+]a���vh'��#??-I�. �^v8�ÃV�� ̻��"�p˛7��X��������I��oX���#��K��|a+���5�#B��sR@HA��[�	���[s��>�� Ԯ��ka�2y{��q��X(����������B�NI09Ͷup��<��s!it�r.�A%���8��]Y�֭w��&�Z�B��@W�1׉�=B�<��e���\��O���'2��F�&�Ns�mݥ���ޤt���#�?�^�����d�ZI~���)~������܃���<9�w��gĭc�l�Q�>𱐨�A�w�ay?W[�����z��DY�.d��Q�Ǝ��X̯mp���p.Yq��>'��r�e��0@�v����`��yƵ�-A
d R.D��h{�p,�u4:hNx��]��Q�2����}1����.���@U�*��[����^���X�>i�bW�4�"dV�n�Gj�;{������H�,����2a��V�/1���?ㄚ��8���kJq��������<JIݢi�d��ȉ�C����d����6�����[.�W��6�k���1��!i푖��6�i��ֵ'�z	<ׯ�)30o�:�>�4h~�0�8��L�ut��޵��`v|��a�)�ߒ[3�]V��c�:�l���n���J�c;���<4�������e�%@5v>�=�-Iw���#�
��@!�a͋��q�Jҳ82RJ��7U�~�2	��&p���S�0��X�:�]y1��1���y�X�k��af�h`��z�%XƗ ���CӺ���D���a{Z�N'GD���{@��'�y��;+W�@�;���N"Q4-Q�L�̑};0!��_���-9�BΥ�&�6��Q���緇��ps_ʥ��j?�.���w=��d���b�	J�2VV:���og���3�Hۜ��尵�n�=��M'WiV������<0����/t�E-"�P�P�YXg���O�9�/~� �� `��8SX�5t�"���� �؜�M�+
a$Ez�tKo�s(�sdq�/�ےq٬���n�{�y��� Q�k���&�ҿ8�uI�����ng���~�pg �V\��[�=e�*���4��7�b�V*?J&�3c�_���U��a�8M��y�K��}GD?v�M�A�, �x0��;&ޤA+v�f1�=p����}���{�>����H����=i��S#�/�~[��eM���#H�J4�6��Z�AoQlP�$�0��hV_�H7���]!�8��I[�9��BB�o8�U8S��a[�`��]���n���y�%>���L�Lw*ʗ����.R�O?�@Ҡ�f/'�j�'�$L�G��EAnuXv���[��	�B��v�a��1E��S�Ӑ�;N��"����"b�����ۗ�����y���������(��Aw�Q�8��G��~X��1�1�d�Ek��#?�.d�'b	���䘗���7�ܣ����'܍���\�[):F��p�c�,�i�z�h�vO�S��?ʔ6�.$a9U�G��Ҧ�W�K���a�^�{����}mk��+P�EM2u�|
�`�n��+n�r#2�ۂ�D��w�Ng�tw��7O&^|�`��P�oTN�1К����)G�MR�!)Nb���z��bc��ͅ�nA[q�1I���_sK�S���,F�lm[-�z�������w#�j�����}M�ڽ"�]��䬕�`�Ӡ�}�7p���t���&�+�0>���;��N�`��[E�N�U7�Si�1�C��ih��;�,ݒL�?��
:�����km�!+���֍��?躕��?� ,�֋H��} oj��$|3���W��'�L�g��	@����d���y�7��Sˠ�#�U�xc.�)`�*c�H3��i].5��[���}����
@�ʏ��R�w@�h��Y�ސ�f��؄�68g���Q#bI¤H�(=1�X*�{�N����菙��8{�@�?�Kx�b�В�e�1ޅ��\S�͈ �PJ�������k�%�֜^�o{�(/W�_� O&��
�d�z�9��f�:��d���k�Fy�JL��qD���.����e�(>c���G2w�p�� f����f�'�r��>:UUA�g�Bmg��?�QJ�M�z�p�<R��_��� E�!C>sR�6��]��緂�+)�e����R�c�m��i<��7g�A��u�oA�pH���Wv;h�N��2����5QD/85��9���y�>�8�K���_�d��9O�I���=v��u��K���
r��x��L��[�I=^i	;k}�$�yT�����0u ����i�g5_���n���oU8���vA���}��+�1v��8�>x��!�
��B	�0%�E������'��9E�klG�ǜ�q�QI�����@��\=z��w�z��	�:��U�:�$���u��X�N�����Y}�u���0:����=L��L��(����ףo�6O�|C��<�#���ū%���˛ب��M���;��V�ד s��a�R����>���tށ��"y��tD'��}!�F�W�v���]��\���9�`&(�/�w�]���>���	�k?�|��aԛ%r��Cr��䵄��8B����N��M��$Һ( D`D[yJ�MZ��L{��J�	�u�nɼ�3uk�o�;�*�ʡuأp�4�r�@��`�}$0V�N����[I��,zR<�g���1YR���w��9�ASWߚ`��	l"�ԙyd��.W�7�9N_Tc�E�X�W���N���ϑ�8���s]� TD$��fp�~��/�W%&�na����n.�f`\M�G<�����L��z�mU
���p�A��0�w�U$z�
y,i�fs7+ڀ��{��|��7�؎�:�1�&��2�5Z�\��;��v��s�@����#�)i�YV���-FOO�R��x\e��N��8��"Mt�ɵc���q���i{�f� 
k\Ֆ&�CWh"=t�g0��}?��;�s��zy�Y�N�ux�M�#b�6Gp �'��A����mаZȉx���N��6E��PD6�hY	��C�a�`�)��3�RIg� =�ez_#���g���p��v���%��cO���.¸������1�/j��]����
f}h���'����nߢށS��-HlIY3��RϷf��c�r��\C�r���yCA��ؠT�v�y*���W�ś�^�$�p��%���}�4���V�	
�!%�&�ep%����K�(�ł�:����D�B�U��1���o`��W��N;��Q1�|�,�۬�Z1��Fz�j������WV?ԕ��T`���ۊY�h���e�$j\�Eu`~Ÿ�,v��g��Bd号�+#�	��i�`�9����C �J��M�SFqˠu�6�"mb�/_�15���t�Կ�Z���V�r���f�lXxO� J\�Sϯn��`	�J����ˠ�O����P�o,hx'��*�U�g�h�jaG����@�p�`@wD`_f��*bCr:<�-��f����;�����U�͟e�m�#����S@f2I�Fh.�	�3��ve>1H�[�a�:,k��}��v&d�9e��ݫs�L��`iȞ���
�(ۇ���6*+x+)�V����b@T��F�j��1�Zy���UZ�W�}��O��
�%1��ͥ?;�l�6@{ߒ{z��I0.��Z��w����x������iX����u���(\8� >{��[V��J:k��*��\�V7U+�H��q�4�ʐ�{�'����gIF����im�x!��M0>{01g}��M8[�b��q
�фH�f�Y�u٭6��8��x�[�d�<��qO���E<=]����:ߌ���Y�y	]P�S"~��ʹS�l��t|��.����C(��F��f���ӼY4�$� �g۴"�G��pr�1�0���$qR�4vE���S���լ 3$l~�g-Z�^���;69�9_F`pp�!2}u6¼9�R����Z�ݝ�!����G���eh�tB��7q�V���
]}ř��e�Y$�vT��r�ގ�Zړ,6�Z�ا!#C��tr)q�-����}�=_ìР���
q�3�@
��EM����C��DT��x�\WMI��<�:�~�О�X1��g�ʫV�ޛ=d�K8Oe��8����ͩA��I�O���z�=py �����vϓ��E�w7+�ij��(��.��X5���j�6�|�� �+]�Ķ�K�ϟ��� �O�p�#Wn�QL:����_��M��0c}ޘ\�[�-��-q�c�1�i�J�vd;9:FMIoU!��T�c�G�FrM���{�+��IdiEU8.ǡ�~�V��Q���Z���Hk����_O�� �u�o���Wc�$����:�q���{�8{��w1��#��_W�z�t߸��Oo��*����a�����C�"O�m�C����3/��1��ɝ�^���?�-4;��_-�Y߀I�xm#�ZO���G7ʹ� �Cz���U�$"C�2���>�)�����9:&��g�蕉'����K�R����ʰ$�� �ȧC�GX��ul%�S( 4*ܖ�P)^�䍼�f�H~/YՓ:'?׆GAY�<A0�ج�Y�P=���#�ȳ��E�]lL����I���DAg�)�f!���%�U�����t�b��a�&�k:�ɟT#�����%t�0+���fM9�u#p���K�q�w�B�Q�~QƐAW~ޙ���ܬ�`mcM�N&G���=n>c�f�ߊ�Q
,����e�C]W�[��R5�3����b�4�X��T_����߅̙"����y�i��u\ׂP��B(�ȸ"=��:{��2C2��͈�����ي����E�/$C���%��nh��W?u߷��r�E��/�NT���:a9ࠫ����5��ؗu b�N���"��-F(yxS�:�cOWu��~��ZK��m;�:��b�/W�h����\��ҭd@���^^­�3ox��v���̢.�{�D�!|`���m��)��q/n��4��6:o�yq�ה� �pV6��Gp�n^�+��c9$�F�?x� �}����/� c����6�<Pma�Ի�I���˕[�<x����Pr'���<3�^�Y��+�ɠ0���I���e5H7�aM`/Xߣ���o�eD\^��ָ�L���OXOy�P��� �J\�8@��x������
����Q&�o��bQH><9^�����u�(| �86*�2>����ᴵ%��L�>ǋP���������w�P1CkK��Kqk��z���S˷�kR*ʫ/]`�A�I�l:ʌ�栓�t0��`�<�7J�#��RD���v������~�<��;�vs��4���1��E�Jl��ɷ�?-/TP~us) ��k�9'[�ݶLW�h��Xq=85�lǐ&=zI�2�V¡[���IQ~��Ŝ��䆭\c��0-���˥�^C�n5T
�'~poSs}��A2ܼ���z��M%��6u�"�ѳ���}"GN��p����A:,�-R�"��kN���ki�k)�*�L!����OO�L`4��\G����O��Y�5���.�HчB�ә�(��n#l
��S
ﮞY#q��e��>�{�
�t �*�4;�T��� m�i��m�ZW�q/;��&2��h�������VN�M��.<��r�O���<攍/^�L�7�� ��@K�i:\�Cq
$�`ێ����\��*}?��RϤ[Ӥ[����;��sԞݦ!�/P�H��D;ժ��*��]Ŗ2��٣��3�ߛx�qr�R�n`-9.��亲�=I2:#h��`���֗
S	�[�2����߈g��*.�wQ���
2���0��c^�0�	�O�Y��QW�E��$�_����tH����Y`��򜍘��*�ያ��QIJ���E)����ֽ��D�>>�KYS�zǔ(�4j��|��[r���/=mV��Uh	����rr��FC=�{�=���%��35+;"O�w��]�[ ��C�eʹ�X�T+�s�:$���c�e2�i����&c��a꺺u���)H���kC��8�>���'��m*8*�����xh�(�3�VɄ<���܂5�U%�P���;��eI?(�GD��c�Ŝ�h �ROah2�zӆ��W��ൔq�)����Þٴ^��P��M�����yƙ�\l�#]�'�I�҉�y�P������I�&��Mz,)��È1����	Bv����"Ab5$(��\8�%�(���'�Pi�khb?���h�e��������~�����;�^��+�� ?�G[�(^�1��#��	��YP-h�IB��=�F�g�$�&X�^_�1��a�#���7��W�{ނ=	WS�Jܰ���s��m����40\e6����,�:|��xn�I���5��qf��n^��{��Q�������3\˜��P����`B/[������w,<�W��nŉR�\N3�70��xʙ�0{���������B�E�t`g#:I4;R[�Ʈȏ��~i�n\��' ���� t�5��|+߷t"Q`n�"����F�BreX�R���b��sAK˭�ɰ9�!�r�Y� �}�;��o�Q�_� ]H��P�gG�QlUm2W�R2oGt�핸bCM���u��Q�<I�4������f&J��e|Ӻ��c���w�F�xN(�js$f�:~�G�]U�K�1Xp�Ž��C���4p[<�X�?&U�5�ً&�;̈́Y,A�D�����0�z8����ܢ2��%,��������Q�n��&Y<7"����88E"VOɛ� �S)"P**�N;bʿ��_1�.�:���X������-�2=��Y*8���-x�J>��l�@��z�\{]U�hq-~Hi�C[��>�a�*�X��P� t�d���:&�<]^yC(<'|��v]�Tɉװ�Z'���6�����0d�b���E�iŉ��FȖ?yt��LI�Vڂ��ϡ�{��hQ��
�Z34��Vɍa֠��i6S�耡T�ð�+�j�؋�ҟ��^�=y�2���ܩZ��4(�	��z�@R�|J)���u��Q�/�B�x��9�:6���XѲ��r�9��j�����Y���w����S�Ė�|AGU����E��4'�.=�h�LT�i��h����y���<G �����L6���/�Rm0�+�֤������4�sJ+a[�����M"���2p����Y�<��p;�Wu*R���������Lo�vj�m�E�וb����ϭwC��Şo�p���S�t����Y����Z<�p@>?^�T'��m 8�# �x�5�&(��M"��	�<3۰'����A?�X]�m��f ��I)��
#KzL<2S2�-�9ӂ�1��r����"V�����W�ݤ�&Q���m�N=���[g��/����!�k|�!��:��6�pk���x��&vrn���Lt��+8�?���c��v�0��p`����''��[�MU40�Ū/="a�#O$���8��0���S�i�A:=����x�2�����D�J���	t� ��G�E�uw�%�ɇz�}�h�r�*׽� Q���6l���.9��5��s^���w.wYe���;`��2e�v���]�9��R����;�ԣ#̋�{١���#�g!��19~�Ӷ�v�̑ޯn;��~Y�f��B�w��^�jCۚ�iݠ���tj?��b1�ʻ�G���|��|'�i�C�ay3t�� ��(NvF��N���u^C|Du=C{�0a����:x|u�?"Հ�.?�����l��gb@�{����iN�k �7��ty���0`F�b����d;:�ɨ�C�T���!����T��>�yw8��P�KN���W��haa�5�v�8&*\�8?�UE.];��ycz��Jˠ���7�ZU�㬇��&����Y}^G΃/��"tf��3J��	�5�s6h] �v�4;4� {؈�-�%�ڛR�f}0�S���4S��lm�S�:�>�� �� �������$�C��w#0�h����-����J]nq��*�w��v�#uy��	cV�ƣ� �:��WT�E���|̠#��_}m�8��g"�Yr\���K�&6����S�s�}���Jr𮫣�K;�L���^8uQ�AIXUɓ�)�P�={d)�Ӊ�H�#e�2�5��S�4:,݊+�(��C�O�"z;�W�&P����6+뎚��ff6`�Y��#̟Ar�zV=�Ŋ�w�`��q{x��J��Q���=K��yǼG�^�;!M�����ݍ�u��7]�N�X�c04뺔��_ʴF%��=g#:�:hF�|��[�;iO�A�Z���+QB�)����Wጊèw�T�^�g�vʟG
nӼl]�����xʓI�`�t�>E��dy�*�.F4��J��prI���T���n5 �h���}ERHa�;�+o��2/'v���?�<��ؽl�-O����AI�cIs��$��$��R��y#���fVK
j��0u������$�S'oM蛴�xܖ��9�v�R?�2I�qj��:��~��ocQ�~O/I������L�#'��f��}zh���'/"����-u�?�:���Ē�
�z��J����{"ì�}/?~�kd3����JH�ڛ�zJ�I ��?Kc��5��FP��*߄n�{֟��UQ�l�n�	��{o�����1��r�n��M�EIֽ�]z6�ѕ?X�o2��˖�^���qB5S�'AeBw����]�eդT�0�'�!.?�CK��@@���_�r�m��m�M��{�U�aHef�y�B%�O�d��x�����2K���x�	|Yl��+e��H�~���bZi���V>>��ׄ��b<��
�ÿ����M(�\;Իqb&�];���5D3RϪ�O$p�%U�is�rswû3�"zE� 
�����5j����.�vP�9�)׃ܚ(�sI�P��_m\w�4���tjޒ�����B�maU7N쎴-��oxjW� ���u���U��8O�և�3p0����!�ܻ~;�ʏ�  �&�d�,<�T��Y)�1�0v�G���4j�p�G��?���1�`ۆ���y�Zzv��B��I���S-rܧ��I�#��#ec)[��{����n찼ĵX���"z����wԓ��<7[%�Ա�%O4re(]ٵvvx�~���i���T~<El�c����G+���3t䠂����Y��g�Lw:�i��k�f���H����v��JH�r~���E�QM5�+f؁PEs��5�U��^n�핅��v+~
H��K�y�"�"��#bC���)?��e
�u���:����I`�B��{�>���=56u��j�e��:�����eg�+z;�i��)kE��+ʅ0��GP��T�y)U��A/�Z$�'S�C���m�Qx�5ȩ�g�zH�(�b��MU���3���@�#�n�.T/yh��s%��T���l�8���I�;q��bS#۳������ �I�/e+Z��s'��4���Ţ�"��\�/��w^�����&'D��Ķ�� P�4i�4��fy�fefC z�nM����_�V~�rIJ`�� ��c>�'`��O*�;R��/L�j.�<�-�dU�+/� �f]y��Z�e;��\M#���I6�� ������@��.���5�(�#��"Қ���C�%�Ӎo�����	G^@����Y~�F�7��o��ـ���2�P�MQp8��~�����'�%�������+ji5ɻ���?�t��l�|C�w�ۗ�7pӼU�[ �i/�+�;TW����W��]1yh&� c����=CӒ9=D��2N@��#K�k%E�B�h�r/b֦�E����o>�2,m�J���5[%U�R�����Jt����wB��R��Q07�	�V��x�*7����6�������Ζ�*��(�q��L�^�̵ l��Aܐ2���n�'��1[@��Ƨ�X@1"��נ�_�T���6,?Z*y2��Ӽ��w���	�'�m#�a�[�����l��Cj�>ެ��+4�H"H��]�**�7��*�pU�?��eh����\Rl~�_ͷs�Ttx9���|!��ZyjdK�r?.Z9?�ڹ)P�M�z��.�$왥̒��_׃R��N	4��݂��5A���N�M��@ꎌ��吰��F���{ՅcV�3�dl�/kI����[�6v9-����Lm���:����J�Y2�b���R~�-s�"���N����٢�D\Gk�H���$�јɳ�=��J�&�}8~�vH�I�}���̔�w��7z�&�^��=������Ÿlv���P�k�0Y��o���gG�4u�|>��mkzF���9rz�uf�R��>7�;����=N��*���u���y��.�5	�nz� Q?=H�̦�,l4���, V���'�QN9&ĢT� �jJ�Ս��O��A6PZ!+�	�Ԗ�>M�h�K�b�]X
�z�g�G�=�cד	�$,�4:E�qI�2gY�����eA袚'�}e����%��1ߊ���,��	H�8��R�Ak�C�Oh�H�Zm����� ��.e��t��	����Y1�7�B�B�>t��l��~�\��� ��r�v�Ov�e��%vQ�x�m�

O@/M����^��v�1��o��+`!'�W��j�w�N��$�:����
(/����,6gYߣK(�O8�Rtbe�;_�%P�3�˛�W��\��|�tp�������h�z]�]r�̌W/�_���M
����"���=�Vkk��s��x��"(�8�ӊ��eW81݆�&�UI��ڨ�9\2=����Y�8���M�iFH��ٮ�Ox4p��e�?�1rc�x�EF�]�e�ӻɐ��v��d�qc�8R�Dz��/�#/�w圄�����J�����<R�o H:,�`����!�����V#��؍�G�!/�4 �u��*�w���=6H�3��!�L`"W�IH������jS}LA��=�(c\��o�N!�8ߔܷZ���RUӚN/(KǯBQ]`�,h��yy�j.��М�x��[0���[;�s�I�ASU��Y�#��9r[|�G�z���d���w�C,u����B�:���8p�����1�\���8����E�`=�`��D%`Ae{oTF6���P,���+�>��t�t3�ƂN��umf��Ū2���Ujݢ��T��+����־�:R�fs��5B!��Aa[��{S&:��7<d��=0��w ���(�ʱ���42Ck|\[gs�J_I1Q�V���h�xE������a/Q/��r8tO�:�^38�.c̄�*O���'1����sp��n�ӕ2-\TfC�ظ*u��g��K���|~�N(��o��{0t�B�}�G�		�/����jym�/��0����,��\Y^a����[��5��ݶ+@^R`]�
G"'!"
���?6Ռٖؗ_&NL�*���� E�z>E�!��x�����DW��Շ.�>z����,�M���a*zE詸&�$���g�d?���;�ki�� ��:��W�=���_��Dh�2u���	��a��vtC�9O���5�����\�5,W�]��
d��(����mY'��𣉱��;�K�D����u���!Yv{�gm�:��z�*0���+�KR����PU�	���Ҋ~�Q %��=��͍��w�?m��S�ʆ���;�YgܷDg"㩍�-���k�L��;K��g�FǀM���f�Q���6�4_��*6����5�x\'*������Pr�t��B�<%
YG�Z�d�>�ѫ\��^}]��q��0�
��@��ψ�R~M����ѐ��_�������<�#�ʱ������K\�QA���17a���)��1���MSF2I�*��u�����ߦN����~đ���<�{���"��ɍ��:R�nO�m�� K��f]fw�lzib�����O��`z���hM3|�SM�+g�|����%g�š�����ES��EW6� 0-v�TYH(),U�3����Z2��c6�Hl������#�͑���ob<�m�C��os��H��̲םa��n"|�fk�8;j�ыN�E'5�OoXK�v���8��g���Fv��H	��Н�,9�R���V}K[F��!��u�rd��,)[֚�y����?�,u�|/����c�P����!�Z��V�,�$��@�X��������G�.�h�kg	j8���F�{���y�b:���0��t���
�p��/`�$
�H3��C^3����M�\��[�̷��n@K�4�B����H��ԇ|�;.Bn⤐R>i��N=��`&[��5�ю�t�I�$��z)A.�pR���0^��X�(�hN&ΈB�.�Vȣ�n�~C��y�`'��d"����nU+%,b&�z?��G����`��O7_pREz��m̬�v��~�
2�^]�����1Vg@}�<�5�����'���u��Fl��P�`���)���#�����WX���B������q7��� <�&�z�)��O�F���+���E�ZV9NG�	U�Է�����A�T�'n�x/zK�e����22Rh�}ẵ�^�_D���)-�; �]޻-9���__���)x9!P�K�)F�Fa�<�+�ޙ��
M!����pO�:�"��sf@L��7�w�ĀKv�׷�;�f 2��)Ȃ�ּ��ۦ��∡�5Y�p�����,̲�-��AD��������\_�T���3��ŬT/l�\�S �mP�;zȟR�V�]�Z���b4[ z���r�`�����x�m�d̈́��|�&����m�A��"]q���i�裠&�+w�A������q�s�
�-�}�]�,/�Ӯ�ɫAے)xpZ5$y�3@�Hd�ws̢�f�� f�5��ͽ؏�ݐ`}C�J�D�qA���My+��*�3ku�~y���h�bB���%Ȥ��Xc�/ ��VVR��Q;�Ua�*��������ʦ
���7��7.k�4׳��~�0��ČE勴u ���|_�yڢ���ײK�[�v Q�-��Mu�@h"Y��c����x���>�b�w�T��fb�dn�Z�̶(������RîA�V݀���/�������ȩ̧j�<#x��X��1��`��}P�x1�Lu���0���nk��T�L!�<V`���z�Z��ʉ�,W��C<��I�N�����E�u$B������n�B�$��pM"�6E���:k�ɴă� `��e&��,�S~�4������Oy��a�y'�w��	�JW�ܥ�IدQ�H��=�g��<�؈9Ǭ$�����FgG��DW�(H��I�z6�N?�{���B��y=l�s�7 [�2����4Je~5���[2|���|� #�Z����W7��P��%\�Sp��C�؉1 A��'
+����0�=��L���ˉ�B��rf��-��f?�����$��_�6RHkH�l�叟U������>3��%#Xx;�VVV�V�vh>�~�<�e�h#@��kt��&������b�E�r�R�#���;�6j�FwZ��Q�������w3�$R-}"{qo���ڐ䉊�X&G�r�l��)H�	�9����N�v8��Yn�I����H�����d����p%��Ze ����}�;��\zY����U�ϖ�C���-T{>jSR^��$=^��s���/`��L��s���/W�>a��-����RĈ�(w���%G�wo]&X��I�f��/��:�"���,L{��J>��'�ԡ��nw}�PJ�>���m�b��g��cl	�H��v=D��ax�S���jFӒ�K-~�M���ˑ�M�}���M���LNT��Uײ��V�	�ǡ�]��gY�|�F(�Vy>ř.�z"��/�Z��Y��d�h��b��v�ܸ������s�ɋ���L&R��o�,JA*w�L�FP��v\��kO�!^2�ʤ����>u�R��𔅕��؛�	�q_����u��h�'y?���)ka�v�J�؆B�5t��IG��QN:8�wlۋ�:<$o��r�����/�p�8�(�'� z��B����� Nk��)�(�F|�w+�Ӏ��c��B쪥����^[vz�fA^�A�l6���+�ɾgh&����g��U�������a)B+�Uf��fxil�+϶��	"#�=�|��:s�ÿ6��Q�����m$2/qI��O������tJ�]\5R��n��
��s)v�Y�2��+MՏ��w�Ip��*�dS%�)x��jO%ʠ��L��c�lG��
Bl�0�IWE��?d+�W�p+��1�^�'|�؞]��x���kƊ^�(�N�s�L������8ntD4
�O�U��\��e_P���z��ȝo�{�$�9��8�۶V�U@.�(��TpF�,Ğ��ŉN~���%�8�a��G������퓊мɕ8
A�}��kq�}�����_rʗ`���9QxF���!�p��V�/B�O���"�`�En۰x�{�� ����$
U
��(X����AD��2.LQ��ʠ��r�S�l9�"�y-�޴�p�'R�θ)&΂�a�C-R'=�d͵"˦�H)<���X8��|r�3K6M\_���v�k/��~����N^$���i�V���Ȫ��Kb�8~'?	WS��\5��Boy'�揌�}�#��Bҙx��W�l7ݙ�y}��
�a�}���h�N���aҒdA��XÇ:�{�ܳ��n��Q�͂`�+T�ᴩc�� �=��G9��Z�h��?��td�E�X��V���xa@%]z`>%���8`O��0��@F)�:hk�|E҈ ��b"&�5����c�S�?�
,�_1�����ϓ|���2ђA�Rd��z�>O��k������.��s_	��Vi�0����3�a#�(�h�:��2�	����\��]� �ٝ�4���揱��<\�o�ݙ�1m�����.p�Vt�������Ǔ�Z�NS�h���%������d��$��?A5bBfa�,�sܔ��o)�F\��6��Ć�����X�1DbH��A
JbXevP��릙h��-���?W�kَ1Q<$N���4/,W�z��7�x�[�}��1�ځ���(�b�(	�l�ND	�	�b�������S�&��*'�b�pM�9Be,��L#���VeC1>�01�8��H`0Y����ah���JQ5��`1��SJ�aö]a����9C\Q@'�pWj� �I�����U�h`}�j�qU�""�z�P*H�)%jk����~$׼��E?OsC��Ã�aqe��+!�wX�Q�Dk��Q�_2�rٔ*C�T:�hd`�o����e����D�z�%w3�J���05�H!Y�"��74�z��S�ʢR-��1h7�0V�%��㼁,K�nU{ڲ�fR��_!C�]�	�����
cpmCreP���t>�#�Y��
ov5�0���M��K��z�;|4��Kδ�}ۇN�N�n/*<���܍��ٴں�)b5�=� qeE��-60�ۇ�\������d�D��Q����ͤ���q��rIM��첵�s�_Z,]Rb.M�|ؚ��c�	�":��L*@Ri1Q f�	3�n���WAY.���%��w3:�~� �����Ň_��؂�)�
�xsqȜp=���I��|I�0b�A��e�@[���3ǢH�M7���Ch�BjJ3�}7P��b��b�};�J��h���[�b8m�����̖��}z�?b�Q3a6��Z�	����V���p`���?���񲏨N�ַ��$P
�չ$��$������,m���;��/��V[��>.Q��+U�՟x�
�#6rf�4b�qJlxl8a���G=�$^#ا�76��=j.�̮ږ��o	��(4��{{�7��N	��bÉ���k9��T'���q��A Q�RJ2�L���_���TG��S���/������ҫꎻ)p��7��μ��v��&�d��qW����������g���p�in$*��}[�D+~pmK�����:�j�r��Vׂh����iZ�Y|e�&m����ǧ_����axgd7�+�$=J���j>�x!\�~�Lry]N����kRcTϐ�QTl3V� ����X;>v#��jJ:K�'�a6^<����O��ɷ�6�%\���$�5�]]�H��Ev�z����RC(�J�;���95R��.Y��;�3�~�lQA��n0�P%��A�D����k�R��?�P]�/�&H|�D>��ٝc��iA��p�L}΁��#�u	���A{�:Y`��������5q*?'jG8��e!�n�"�n�k��v���Ф��>�t���H���>1�����T����
?g�z�3�$4�$J��hR/�G����q�V��PTD6��Q�l��_`��j��&=�>��C �NG��(�s����/H����&{��)ygBX��m[���2W^c�h|irs?�+�N��lE��ɮa"�=�9���D/�cSښ���S?q��s� �F�&�*��:��\`ŷ��Sedwd�/uj�S���}���&�-*����k�@�mu>��&��g[�݋ғЭ�y�ƶ�cԉ�f����FG�fV����fY��D��,/�{�0������I�-u�^��oP��\j�<�
��"_rX��t���>����1V�8�$�����mhی�Q	_����х1P���x���HM���.{�����r̕"T�#2�iO�H�p�`��ќ�4�r'l�{䫴�l��,�R&r ����֙��Ø}������)�-B���g���'+mo�r��@����;��bbwˮp�7�恿�[1@Ê[�<)�ja$�dQI�2�;@�m�NP��5/�e`���		&:+��� xW�2U�2&��;� ���:��7 2B(l����)��I�÷�ד���Lݹg���WIv���k4dd�I�ŦA�� ������]�OL0�,��j�y��ht� i-�H� H��My��N�2���L�8�~\�'}o���⋬&k��s�lÖ�(����2F�EC��W0�z���:̳���΍��R�
���YL]V�e�ې�6J�]��=qO��ᢌv�&��,��$^j�����-2qK��"-�m�3Ms�V]����I�2�j��iQ	-�բG8��>��o!����ʨx�����.]���R��DC���|l�:��t��Ѹd /Y�Hq����vHG�s龐9r�Z�5�}������E�&���\wM���ڸ�'����B�#�a K���W�q{�x��t���S���v_&�蒳q���
U�3X%C��	M�b�vKu��T'�W�$_炍S�(dcv�B���p�ԕ^����í����akK�Z����ѣf�:}���P��T���f��_T�5:!�����T���]BfJ��Pwg�8T�mxA=,!��-���hC\�����vv!�N'Q���}�d�$�)��$áZ�DTK��u'[\}�t��t���C����QJ����u�^�3R<��f|b�/��:}�U�i�i+RM����ӆ�h��|���<@b"��/�Q�d[�(h��-�*H�Mb�����*��o+U���;{-�e��8�x?F�qfv��
�ģ�L� �;'�}��{��8����~J瓞�4^��� �o
� ߇��`�>u{߫�K��b!�Ĵ��9]�פ%�[��H��̴��w�A���]HӇYE���ͬbخa���C�Awf�x����❹��{n���!�С.1r;��,��L���Ҍ#�gƴ�@	&"�[(��@}Q?��R�"EN���XeVh�ך���F�1�L~\kt�ƽ���78^$��X� �	��)~*��r��5�Tm���xO�����`2o~�L�{��k�kP%k�ԧ&v�UBd�Aǈy6ek�Y;�}���|�hr�oK6ȳ�Q��PW��+m��c�jֿBk|A�Z�H�`�9#!���(��% ��J�B+�nnb���RV-��O�7�5QjzQ<�'g��_��} EM0�_=�Z�}�yp��Ɣ�	7�)I�`����&�rGLi�����ԭ��AoQ0������ǲ�m ���8FQD ��>s@���a��{�s���2���2V�*�0���4�b/���7w���"ti����\��A����쇨��}Q��h�1{J�j�p�yi�%´��%�_aF�瓧�ASyEm>bVw��%4���+�8i
�\��TR�+��ƙ�@�?b�v�v�=��#;�u1�mju��P��?�E�2�|�O�#0pL��N1�y�
�P+�-��+����݂&oͥ@˕z��UN曀��=�}3:�jpL�d���mª���H��8�D���\0X�_a?t<.�1��폆(��)��	�P���_Գq�9T��C�ԏ� �a�Ѥ|�oA���^���2��I�a]������ݺO����q�쩅����:�r�q�h�̚�sW	�^:���-0�41�G�Ú˦�P�q��p)QGαI�Q�|}w)�v�L���?������zr�wP#��d�L�Yr0��y�F�����y?-L��)\��@��ǥ
��p�%�'8��z"nn�*v΁<���~�!�T2�P���oD����Ֆ�82��z�(3� ���=y���nɼS`7�:hR߿7]����j�|c'Ï22��C�%+Z�]�F�Gd�H�Ql.��_��?����}޴
�}�������u�р�h�!2���>ɼ�(��=���g5�n^F���L#�l�%x�Ԟ�^I
�x��\�ڽ��e��^[�)gZ5��jِ�V\���!ycƮ(�}twHckg�D�A�=	��;�hL�{��#�b7����œ����Bdn�է�[��,-����"Z��D+�e��xϭW�9�+�F��/W3H>�oJ�֒�m�~x>j�7X�?�-qU�b���)�Fb��IX�=�@��eՉ��:aҡ����[z)��Is3S}�F뛐�H��S��*�R>;�P���ٟg�*ۖ	3Q��9p�/�!i}�����}�#<���t>#?�j6Yg���6�g/z��g�t�W1�ū���^$�ݬN�J�똘n8�u����Hx�|���l��#�@����p��I=�4�H/^�(� �� 	�=`���p�����*³4�*���@�� ��]S�^A��j
���)Y��MSQ֟ujS���G�i��0f#.N����C��OB@�V5�~r�Qm��\;_��PB�D�*�=�w�����|�(t8�m.LI��MJe��֮�Oy˥�8V5���/H�N�y�s(hk301���:�z��{ %�{)���á��,l<�RCխAàWiC���on��݂4��O-�5�̥+y�Y4_���2{��t6�B��>Gv綽
�7D;&1X��r���N�
�2�����!U�\�z^-?��8X8wМ��TW"�F�a�FxH����>�u����k���K% _�g��]�9��)E �#h\�?ZT ���4�����2�z��V�z;�r��V�b,ӥ �C;?����!#�Tڵ��J��l��5L�>��Q珸Sf��X!N��Q���t�\s~���F
�l�&�A���X6�=���x��C3��/����A�F�]F5�P�sMR� \^��D�z�(�\�\��?
��!���D�ǃ7���J<�f Էs�y������ݿ�^I/�͊b����.����a�x!G��=����
3���(9����{�D��^3\�^��-w�4�i��Կ��8�  _�9-�tn�|巔��5�2��P��C ��dS�I*wh�u?�B��n
�+��qFd�n��%�e�egh�����KH�qV&V��i��ڲ��%X����ʎ���U�K���y��(7𢰾���.�iw�슏������q����\d$�З�H�)�0�F�n$�Z��S���)��s$�9�IJO]/�=�~��1�Z��@�gƉ�_!`1�c��
���`�<�3����N=�����s,a�.��G��I-E+�����ғ/�����H�s!��8��g/��|�y.z��lT�O�RF��#�W���%��7f��ۭ�&�!�4e�P[�ǯ��0��[�܍��u��h�P�������w�����,dM���P\�|Topđ���Jk��N����˷S��A���QkOs�L��wr��=�BN����D�5�jD�v�i�|�$UѻP��q��n!&
�\�-�|������_AlWB��x�d�1��_���R���Fkk�SG����#�~�%��gA,�b;B{���f0���D�@����B�*�4~��_Ǐ虼�yWw��+�����?.���
�loQ! 
���S��)��G> i��q @�R��a��ra�n��M����
�6N�$�3�n��$��M![B��n��u�,��!<ʷ�|��9��A�J�vGq!?�����J}�_�7�~�$�r��xZcIfB�b�z��i\.%�g�Q�����-3�m,�H���W�4��O'9B�y<D�V��{��LsX,�3"����S��_�i �N[]6Q$�Wuf�7���+���,s�x�b]Z��$V���ik��L��	�� ���T�zot���Z�z/�g9:�~_C;�7�ޣ����"ʡ4˄��h@���$�Aa
���l[���'��[��>�7%t�v��L~��6m]ˇ�?$�U!��J�%�S�0>�pM�O-r�7.�N@�6�<`弯�;�5�#6�8�-UdƇ���j��c��h�r��A��P`#M��v�$����T���{��@�Ù����f%mYK1�%���T��.�º?�����B�CY7I���xɝ��C�F�G�lDho�Ӛ+q��ZH�����-���=tI"�a�H���g`؊ ��M��T1�tF�u6�>t�?�2������i֗����+]چd�ƥ����	.���N� T[!n{&�d�k����wDeH�FMspz�n#'{a�5?�[�ԉD�״�_�O��@��"���S�w^��ߺ���Z٪5K�
'�:��.�����:���' ����j;[�wQ1��4�ʙ^����u_zf�BG�EMȮ������F�K���[U���1��B�Z��ם�JA�pcY��Tʶ�TM�	�PD�(E���CN{+��SC��/h��zhB��6qe�j��D�|WnJ�$ozU�6��Ǻj�j�WM��@�>q��G:���޾�V�˓�'�^���I���KQx���WNa��5��0�ޕ=dë��'�(C�L�,�#��b;C�* �S��xH�/l�����]��~g�B��M�����L�C�r����z�-��N�~����seI���,���M�s������{ �ff���/|��*���fef�q��@��B�"������>t�h1Ϩ�aR�z [XT�2M7���f�;_�C5�n��{����_r_L����J��x������~�0�+���x�bRؖ^W��6*���{"6H��q&u���(��8�i��p�Y��I~#t?��_�?V��}��GAmc|Ѓ�6�ʩ6�iN�� )ti�|W�mF#�]���;J���"��#��Gc
ǽ�/�o5	�8x�P�6O�%�S5B�{��^�0���ѿ�O	�;�"�r���Izܪ�#G����Ƭs���H{{:�,��k(�̾�A��S���s.O\}c7E�r����	���sU����Ҏ�6J|c�r��bN�/�\y�el	�BF�gT'��@e	��OAhC��;��R/��p����[~2H.P��B�3T�7t�l�ߟ{����X����A�oK�r�i�(�����Z/��K�R
���q٤��]j���4�UW#}�"@9Z�yL;�K����R��ѭ֜<��@�W<���+�^�q&=oO��Xx����^\�$)��z^�w��#��a6�^�RV�T#"��׶B��}��K4w�$)����[2�ĕQ6�J�\����Փ�5"e۬M�����W�h'E-h`�G��b���N�z*����+Egt�_�)Q(#N[7%{����*-؈�{��>ׯ����2f%�yuʾ3�̱v"�9Fe���8.L�U��Q�T=1rq����lnq)J��d�	y>�9�8��Ru\4��aԊ,����FPQ31��z���j���r����q픒B/A������Ty!K����./�[��tq�K ô��js67��e���)���V�*���Y�'&vC��٘����k�K�?��6�=��T���r�|$�ݣ�P��e#������ܯR#�%�e<Q�o�4U���;+5�F(O�R.�M��J���7���C͊�D��5">o���D��tDkC��F6�E�+��5`�2+���J�Q��Q��:}F��ӔC����c����=C����^�&�0��j$=v?�a<�	\1�����0�!��.��8D�ӿJ�� �lk).^�:�~�S�`��(�K�l���0�6J�%�H"���S�:ˉ�D�.��/����M�ݢ�M��Y%Y�y�:ҵ�(�x���e������Xט-\����u`Zl�J��3Ce�c���h��g`�J�naAm,#r�"�P�s����)nӷ���:�]6o�&U��y3�wHA��$�>aKM���_.܌9� ����fuU���)�J���ҁ��qi��4�>e�:�.T4���d�ش��M/�Փ34�y�Z)+�[
`�a��sUK�"s�^}�������D�4���5xe�i�����b
@��8Vml,�We{���BeƯ�Q�h����$���*��:$��F}wX(-��ߑD����\>�+i����i����q���*&��ֺ�>y��\#y�~�A�B�C���$�7y������w��	t�5��##��ް\܏��������re��#4eC�_y����� ��B�nK�se�*�dbkŅ�n�`n�6�q����V���ӘX�`a_�����QXKNI���7�۵ronz����rY���'Ĉt���N�/��U�Ns�r������斟��b��4T��;��_��%�b��㪰'����d�J\�0�#�U�^Ʒ�W��bVC�}����nE�Μc�BѲJ�r��m�50��D���z	��Ye#�Ϙ�Η�2	U�-����u?���=s�<���K�dU�S2G��R��d�HYw�,��^ِ.`�X��^=�[(~( p�͚kPhl~�2�Qf�9/�b]�~�>e'G�;��⁠qJB2�����$v��{��=76�*���'xv)j%`ք�&z�{�^�u�^��m�j��,f�H�Y��N�$��6�\@����]��"�D�)�&~�11ϪI�\���1wET�/�c
�Kf��b����N鶹���g�~8�Dfީ
j�%�!�N��g7ȽƖ����T~���jp�ۇ������m�wrph1�L�Ohe1���޸{�˭�;e�]"I��^�������H�
�O(��U��oA�ٲ�@����ߜ��������=i������6<��8{��OP}����R���A�Nޙ9~��%NGϔ�Di1C�<0+�JdSL ψ��w���XWf��ͅfc�I��u(YH!e+��b��΀���=�mml3�X�p�Z
�>�hF��R��iБ�s��G����I(����X��u�=�A[a�k�����R)���=D'��a�@vl"[��YSd��|�c���Ž���y�-0���M���n=A�5���FI��p�7K����pX��Y�t���&��M�Iao�Pެ��bU�]INC!�o ��$:#�ELn�iߔ��v�3�k��"��]��={������c&!B@� A��sمf4�"*Js���T�	_��:�b�Ky���t���W�I���4:����2i,�h�U�qMn���-�z�^u@x��[{=�ű(�ݧsF���r����G���w�R�ۣ������yv�����E���OG����h����Q������T6�;����a�O�`��fڑ������&h�'$�͚�֙����2_Z�x��/<����5m��N�6 ,s��Ҥ����*"d@�s�N�k����q$WfB��ܼ��Ҫa�q\�%�;6�	�/������R@㶆��K�����딝U�#.��jA*� �%�Hg�^�m�S��%�Տ��^*ψ$�Ԛ�'2e��Ԟ���C@p�ҏ1�E�k����Ȃ3��BJv;x����[�)B@����HZ������]phgS�CHzF�)d$��ϻb���uC,���Bf����������u ��L]�o&��tw!�C�q�,v�?%��*����
�=�y�_C��F-{�4%�j��H���S�5�/5�tĐ�_�}/_��M���"R�o���X�K�dҺyH5��ɔN�)C�yL�rb$F�Qs؃U*H*o��c�Q>��?�����K�k�\�g��K���iP��	r������.�0$.�3&��*ttO+7C3���u~{�g~?	�����_.>�郝��E��녂��I:$���-���\P�E�� ��5�\C����9�%�#Y�+������Be�ׯ��uH�PbG���oO(�(ILr���a������1�ha����e������$�)�f�*L'J�	����(Z��0cQ��>'��0B���z�����fT�ߖ!���x��Ҡ�y0o��>Z=���D��䨧�m ��meCDm��6�s�7ȴK0��o�^p`���4Q�Ef��"��9��,��� ������¦Wۖ	L|~�-9Q���Ŭ"^��� ۥh���_��1��2����vu9��\��~RGn�
�c�%ؐ�9?��ic���e2�H��.���T~t���WȺ���#"��D_w�<a>F�����{��h��.��S�5���̎��+�6No.�b)I׽
^�UE��	�IiW��E}jB81s	<)����h�Ib��n{��/�v�q�B:hI��ՠ�,��|����`�)j�s�0T�4Tw�� 4׹���d��*����!��L�=����J^�>>|�-ml���	�8{���7���X��G��H�B5�T�Đ7Xk�$�~�@��9�*=3�zk~����zC����$�
�$�5]ڰ�#D�G*s8 �lVHsQX��F/jX�k"��8L�p𩜳C���n��0O���\��e[���E�/rh�2��$.D�j̼�m�`} �Ȫ�H�����G��B���X[aȪ#��v[o�����ԃ�m�U��������C]rx�9Bu!ʇ��0kv:�J��������]yW��#f/�����	���`���6����}�ц��sI-���WX �a}�֬X\
,U��Ihɗ���j�ؼ���9���J��"5	�����n|��k�V��&�ϔ�U�۴S��%�
gw�X��^Q^'���3����FC�z
�X����Ʉ�g�Ch̜�G(���r9W��h�u�Q�,U��5sޢ��ɢx�w��������$�e-�g(��r�uC�Z,��Q3e��fС�Lq�ˑ�hF6X���z��)ͪ�dR��s�+,�"����'J��e)�$DP,��>{���dʽf�������ߒC��z|J�dEh���|&�S� 2��o0~�h#L*���������,�� +1�I�k���Vu��nׇ{�z��=����1�x��^�W�9��H8	��_�.�z�m� ]��$�m/�Z3-e�*�EHZ�>$�W6�ן�΀*&p2oTkH��rXy.����c�I6� �`�?�$zΚ���ep;�c�{&�<�JP6ӚQ�A�U�8;b��x���#@t�K�����1즫0��=�\.����?loGE�� �{D�+����4(j��#.%L�_IES���[L��ئ�0�]�h�g*�mI毷�S������n��{�Q�.���_~��"��7u�%ͥ�0׌��tda�ǛP^����< [�RmK�qܤ\�5O��UbL��*��
�P���!9���sf�w��$���gV])Ot+�Sr[sL<z��H�/���g�(z�3��<�]Tڭ����hr�O���.��6 \�W*����L&LՓ��r���76#H�\z��i>�͎B6�x�%�����@5�����-�}�5��.�L���Qw]5��/^��Py\�D��Ye4�٠fhf�C�Ds�y�<k��>;���gTB��n֢����jtH��}5�SV�u�D��n���
�:dQ�D����0��.��� �7u��<Tt�K硂��o$�F��8�缻�?�d�Q\��26��Mj��R�	�G�4Hk8��[�q&����땛 vC-���Լ����h\U�<X2����z<�ʂ�1�>�u�ƉK�D`o��5���x�������c(�c^�F0���h�SI�ZdG/oi�\I{<�<tu�.t��@��G�U�EK��4á���N$��x�J���Q{ݬ]uD}YV�8*P3�"�?�ob夆aa	9�aTj�]�%�䐤�t���&~��N������%�=� ����>�G�?5�
q�^��e�nS54]p +��1T�Q��P�*��2����ht�Q���/`N��C��<44�Z^�Z��$2S������qp7�#�<fK�2��W�>��L�E���HV�Kk���B���rS����?e|�9�B╉�p����Pi�J�F��q���|���yÿ�f�k`��� �@�����vJ�d�2��	�x�A�&*3J[w�RGu�X�����Tb7���Ý�ge:���x�J�\M��>?�e�4�0�N�d��S���������m���_��=��~�U���$�vx߫!j=�y?ߵE8q����"��F���8�*�Z(Ojpa�������Ol]��'\��<�lX�kNi憟�O�#�?lۣ����R��ɫo[�v�<�%֩H/oI��Q9<P�z`�5����~t0�(c�E����0m���cA<(p|��>�5D�-Ȗ��R%JG��0�-?˻��b哃�?�` 2y��WQ]�&��w��"��l�/ko��Jm�G�Sʊ6����s!&��	*�j��i�S`\���K^�,�To�����2����j������4V�M��"�e���foܐ��sݑjH��5G�I�꾖�1v�?I�H�] ݚ�]Tt���^�:���B��:P03wr`)�(��cS��?�*JD0��V�%�|8��q0¤"�肪-�8��r-�nb�j6�qG�hP5~	�e�����q;�֍����t��f��k�h��IR;����{�:�V�6]��K:582��)0 }lS�N�x�s�h� ��`�c��bȃ�;��`�m��x6Jw��O&��XtO�#"����|_@�]�C�Y�=��I��G~bȿ�;�ZtzVPJ�,j 6ZcH�̩�q�������u�K�������P�(x�E��6�ڄp�΅:����;�ǵBJAm��Y� ��)dៗ�`�c��1���{�,n��㺋���p���V�L͈Tړ��Gx�#���7p*/�7���!k�N��ϔ��س]~��[�m�:s,���h�2�v&����$�;[��#�CѼ�fÐ�F;�,pn�gf�+�M�O��	s)�d���|���Xc��%�����d����#����h�i�}x ڜ���]��! ���v,CBMl�?�����V�sM�����;�o�+oj�()O.T���:���a[D:>�A��h���绞\� q���p tx��N�Si�P�Y�5�����ڰn�C�[2�N��l�(���-��r�iB @�j�y��8 	F����j�I��	O��hI
Q+m���J|��H?�&g���wO5��ª*�F`d�ud����w���R)]�t×�S�P�����aT��t2�ɟkHwU*��@'ڐ��gB��Yn�o�n��U��`ċih8x�Y~�x��[��������R0��N�g��nTEѦ�?�ob~�bv~����Y�t0�J�K{��ʪex��L��iiv7ETh��;cH�~�HY��Ǧ���w��9��5����׭�o<	��P8Z3��v����?������k��n"!o�𖢙s�j
G�*�^- 3��{�����H��|�=u��{�r�����`�� ��l�DGZ&��&Q
�#j���rO�%[�8��t��׭�9���}�l���j,=:�y����p)���n�����G~��?�J��E��z���?.&�f!���o�i(�T�B����e��x��5'
�B�S1�`�i����m~$�\�^��?�с�� U��P�L���*Q��G)8�a-g���R��#{�ej�M�>�R���L��ٸ�=ݰ�D��=�Z��	���-_2��8b=ǌD��F޹�������UD.��u�a�� -�����E��pU/-��]�F)қZ�饒���3e���EU��=K�h.B́����%U|��
�<q%��8��{-�̐M�F (��/�Q����|�aU����RY9`��o��P�;C�`?Zi�M� �SX>7 ��>�d�Qmu�AWn�q�]����q���=�E����}���\KK��^8ĚD�}����V9����G����)���T��^�sD��u׫H�$�FR��t�zڦ�>�X�ߠ���P(*�M:E;8M4���;��J\7�G���&�����{4����uܝ��Ds�U���y����Se���� Y��ZqH�חX���V�C!mI|]�p��V^�%��=a�jcY� %�5���s����Sq�1�KjY�@�<��o�&l�A@�k��4�n:PB���T[������
I\;|?�9`�#|�o�e�9@9VX�馰����fɸT'W�X|r�5T�Bd��9���&�
D0���K
��l|���j[nI�-�\�2jvp�d�R7߰�c�p��_
Gf��Z�����P�i/wndd�1��ɓYL�ds��Oo�M�Ï�)�9~�tM����v{�DQ�f;�	�,zP*-��KB��j3�;��_�u7D���K��F�@7Ų�����9����V��a��������Rc���r)0�$��݈9�{������[��]��ٖ`���
x�G>����g��k�c��徳ǒ�WE��7�� p�̀�a1R�5��?@F}�8�ڝ��Iw�dHY�Ը��������>��|�c��*���P�=a����a"j�_p��Iݭ-�^:��/h���M��*�@O�/�s��@�{!Ѣ�.L�t�JeT�p�m.�Ikj��4�1����$4h�/�p)�k{�9��~�$�V	dk���TMGaBz���s|�'��l�?�:��4hޥ��T���Me�}�z�F�� ED*4�t7J/�`��v������i�Z��*?��CV=�݉jїcɆB	�uAģŮ33Ŏ�m~��M����{^�����+]�c5@��EQ_h��c6~�b��_�Bay�;4�6�Q�ϜH�c�:��t;�,3�CZ��c蛾b�<���a)�+e�7.�ʥ�1�ll��Z����z�C������S���K��u�Щ'�M�J<.:3��+A/�cOON���iV�]�7qI��zWe~;^&`�ˬ�@m�[�h��a�+r�'�IM�O�C��oD�s&� �I��U��8X��]����3��]�q*)����i�75V��S������z!.����3}z��@���p�'��]�{KN�'	|��>�)��QǺ���W\�lI���{��P�hA�:�d���Ũ�m�p�~�Fqz��מ��N�!��nPu�rzH�
���g�	�+��֝����;n��ꤨ%��n���F9���9l�J��KΖ���w{�8�x�oO��#���5������hc|��~����h:���0���Te�v��U�!�ܠo2���F�(����m� ��>:�~[F����-+v/Ǜ&$þ{�ld��߄3"���p���GP��fvw���܄���=,��(PJ�I,�mu�*8�N����^�
<���Ho}K\��H�4o)��^Ṽ�U	\�j�Q����c[K }t���27�E�F軩$c����5���H���͓y�g<�8Z���k��0�\D���<�O ���9U��Bg�XRDo��Ө|�Uh�E�W����j~��Q:느��H6��y��O�-,�9A��NC�-i�{?�8 ����9�&E�S�ym�h�� ��?�� ��'=�Z���:�Ơ(�M�Zg�ĸk��ZXe��ܘ���^�N���X���7@����_�H��s�fPjf���9҈ V�����|[��>~lZY�˶����x�硻�@�80��M�����~���5�����>���RC)��\��v�����ڳCR<ue⻳O�����t��(gv��o/��U������+�!��bD�a���v�p�z&!lR7���W� eɘRsv
ܙ� N�.�ȥĸ$O.!���PU��慺�Ov������u�G�;�z|m����,���@��v�Jo'����4H�R&k�� ��e�f��t?p��κnU41h*g@"ɶ#�Βk��RjR���Bj��uܬ�Q}˜M�Sq~��}�ؘZ�V15e�
�>�O�g ����՝�:0�#����J�ni�D��0�R~k��Î��r��vG��ρ �KV�r#g��U��[��� ��Q����;�СB/�z���*>+��8)O�Ne�������j�0k�{�}'M2��\�b�D][K�ޝLv>����Z��''W��k�^��z�A8.
�W�mf!�[��S��B��#u�@�%f0"�����)�+�1�[�	�Z���B�؉
�!�o��Ê���go��d@�'���W�]��sp�"w�%��ލq��}�(��>�e����A'��7]{��d4����9�#�Zs���rp���')�eV_�1t�5�=�w]�����`�
��P�.��Bt��IY�$(�h"�6�'0�8`���"Gӓ�19\G<�(*�ۯ1OL�ُ���z���ԎcN��C����d-��h��W�^�"$&�a�vn}֍U:u��m�ut�Dm��W��Hc+(�\fO�����Q�ٿt>JX���<�`Pp̞����&%Sp�W�`�����L��T0!����a�D��[��)?㋮���ڭ� Dՙ�Fh�G�8sPD�"i�ň��	;�ߎ5T��S�ۚ�_�$)�XX���ԕ�
�w��g��N��~���\�S�$�x��,�@M=_K�����Zm���m���V�$�Th��T4�����xo����pS&;D���6�3S��v)�����gL9�|M�>�h��E��$��W���RI��jS�i����:�oh�HP�DNx$3�,ra'۲�=SL�I��=��~��$�W)�Rd &V��ޣ��������C��cC�!��=�3D2�/�����%��F�:����+&��G�`���0Z��'�����?��a���M
&��U�f����=F�#���t��ۛ�I~�3��u_��w
��S`�Р�t�,z$��Y>Q/�7nώ��yC3�`V�9x"��m�ƧҦ)8mve�ޢ�d��p�����n�"�R��*KL�tb��R�B�,��l���-��)����m��n�E�Tn�-uql��s6>�!�c�����@�x����Z���۹@������T�"�b��J���.1@�j�a!��A�8'z�|�,�a�Q�oZ;p�܂�M�q�
J�|i`	����|u ml��2n�^*Xy"`kn����"$l�w �6�tg0��4ER� �ǆTk!A{�@��^�`����s�L�ꋋ�5d�����ǔx�����5yfRK[��m8�+Yo]��W��"a���k��O�x+?r��
_�!ya� l)�zȍ�ߦ|g�A��a��.hW�l�%xD�H�G�J�mĊޙ|��.�\8D�ߺ6�0���������ng^���K��g�}J^W���kc^�uC�^��$��q/"
����[�l,����,HYp�i.�0[��M3�`�.��:�캴D��E��XmaxсP]_��bnc�$*W<pץ|>��T$��	�L���(Űy���=kYHJuRr�����~K�k�"/x�!tn���K��;�yU�vE�G�-�#�T��Պ+�6���Ͼa5|0<�1����T���A�f��k�iPB��u�V��$Ƙ��;kN'ZS"����������"���%��b���Q��nd��2f�%�Ŭ���,�/���<�0ܸ���(�{���ͤ���P�j/�������v�?��g���mUQ:�a�=�8�����pG��A:�&d�xޛ!�7H���}�1�N͔Ƕ��X�������s>��A��~ȨS,��� _Q��u���w����*��3���C���*������	���.@0DO4�8��)K�Ȱ5BIJ��_��=v	n��_b��^"�@Ns�*&H�H�m����\�(G���b�&f>��㟵7�mC�H��؏�h����r5�"E,=���a�S�ޣg?*���B!�væݸ�DbMzW��I_5v@�)ѿ�>=�*�%~���\�����V}����H%yR��%�]c�B��|?�طp�W�J�o� �6ц�3��}}M��H*$�7�Su��p�e������B���y���^�/߂wͩ���a�qk��� V��
<i7��^�:��'�۪�J��H���=t;�1Q;a5i:�tBXAF��d��a1˖���A�k�&���ޅ^DIxŝ�K��Vo1�����J �vp@�5���`�65�O���e����U�J@��=������Y���i��1�Ɨ�y�j�*������
�l�r���1@���������r���(���/_@;�Z��t������~P�����`VU�ZS��u���
~�k�/����a��:��`����������r��e7����Մ"���,G݂`�3��k֢*
����=��y�a#��T�5$V���\-�')#jx&��7kgt��*t��bHx���ǒ9��N�?R���7�����{s�0��ɼ�{t��G%D�C�0��=L�I�����QK�d�Ŕ�Q�CMYsAG�q�Ao	��������e�z��cF{N�&�	�,*$HP�d�}d����.�,7�EL�B?��p�^>=އ�gBZ_=)�Ζ���
�L@��
��� �&�H�Siߥ�G�m�7�O�yQ���1��'	%���w.���.xu����i�fJt6�_�cк��.��iC���e?��a��nN���[�.��Q��K������"u�9|��M
>f�.�����j�z�t)Y��P�z�㡠����ƀ�P�^�&��Q��5Y���ӭEG�ͯ}�0i�T�� �wfE�A�7ˆ����-�-<cK�!�ix\��瞌���R..n)�)��וu����B��D�s�:t��Tg"0�w�Ԁ��T�ZZV�#�eP��d!?8�(��ٻ�iس)�b��c	�wx���-�I�ء�j��<(XR�\�흔�� ���#�Y��9���ʢ6��Z!`��)�:�XҰ�X:����Yw��I�� (��bƁX�~<N�Ŏ�p0��B�07���K��'`��Ʃ}�B^�����9��-���J�5O�=[wo���(�<`L�<��k�|�H`7t�Z�G0 �s�7N|�@�_\0���^���k~?�e-s`r\C;����}���$O��!����V�m���8�Q�a^*~r(%�C��.��$N+�*.�{��E��raJ���)�(�N��W�7�`�u�?R�{��G�c�S��Զ��*�Q�M׵�<4)�m2+$��!݅�^���`ߥ^�rAp���"N�-�
>z����a�	X�P�t���l�0��b�nXM�~�j��9�fj�_�4�EIGra�O�\��[Ս�?���h��M'T,d��2-�X�<�	t�2��+�?���Z�����-Dw�]ʑ�H�Jdûd�����=�|S�ja?�hU�?��8��ڔ�ğ�:�����C�(�x��7�lD-5��ʦu�v����'*��݁ō�O�3WJR����hjƦ�t��x��6'Y8�M��Ed��९�H���x�����.By���\O�����Q��3s�B��No���@e$�ƣ���p��,�٘z9Je_c
 S�(X��{���!$�fۂ��52R4`sn�Zg;�FcǞ��>��#���
���'��O|�*,y�W��fTCvP:�?N*����Qu�}pu#T`�Z�{*Pp�E�NS�幕3_h��|b'��'Q��{��k,��M��gg�y��s�4�'9í{����&���%�|FyE�_�8��w�d��q�Ê�_m�\!0I�:v�\�O7F���+���g_0Dzˬd��9�Ε�C���֥��C�،�1xX�A@��a�0[l����G�7?�RPt��Y}��v�#;k#�Ԣ�D�7���xȱ�34�a~�)d(�#��B����3ZH��7����%�p�?��#����n\4�&�Xk�C�G�,�Oڽ�2庾W�ۑ�#"�f�FE睦;jC[7�����,����`}���^cU�@�� /�򧏈Tܡ��A�յ�Ȝ�t�2�lA�5EO!Q*$L�M����W�U9��Lw���ԙ�1�ɫ��DêZ���u"�nd��T�B�`�!��뢴����(����m�"�V�vuJ@�q,��[rbU��MmHv��!V���#�E�5ރ�)9�<W$�?���W9�,}΋sхJ���lpWEc�u��)��>)�l.�<J��8�K/§�\^ۑ��@N���:�C�<�W��;	�nqxY. j�V&�NjGAby��w��ǥJ6m[f���򇑣y������8�	��7�����z
�8"Z��I�B���gR�#�p'tƝ�	yb>`�m��,�T:�J�f#XD�O�3��'O2��c�y4���G%T��T�wђe��:9o�o���3u�r�������a;�&�ɽ�f>U��\�*���g�T�� �0K���v]D�e�X1Ȩd�j��)ܸ��X�����9�j ��3G����3:g�\?�a�O�4�6�Z�}��o�oE�#4^�ObhCr7����~Tbjjp�U�������Pg�C^uM�o��Һ�h�I�x�ʦ���olzud^ay�M����'�v�~`@���4���r
�ڥy�� "T����G�a�m$�����Q�.Ō>]��!P��z��N�C��	�}��Cۗ��Ъ"�_9Ȩ��:�Lk	+mh�ܒ�7���̊�I4��hhI�_`��?&䶉�l]� ��xɲk���L��iy���ύ�{��DP��F�DM�:�9ɩ��h)���iG����'"hW�ͯ���[Х?�Iݔjum�� BR�O ��>�0/�t�,�f�3��{.�1Z�p�I�9'��r�k�949{�:�H��I&�]��MnFw��҄�v�(��o�<Ԯ"V?����j>���pQ�6%>u�2��Ne`ey���X*��o&� n�>�	y��N�ć��,����h�c��וy�i�^Ӧ^������=���D!��L@�2_��t�ȳ���"����-9�v�[[��w�oT���9�釦��T�¹�\oCa#!��;��=P��wjR�Q���n�S�o�~
�!�qT Au0�ts�q�����1�5؁�;A��	���S�e@!4|�ȡ�?`���se|v���5C��M{Z� p��ِ������B�"�?
R���O�r̴gD��W����[���w^w`���D���[ �Ώ�"��@a��Zd�)�r�^�"%��W�96��К�k��x]!hGAH��sB���3B�0
�ܝ����.y��p�#A4��m�Rc�º0�Q��} ����fcs��F�+��"��'a���@��n�r�XK����?�v27��*�!�i�nu?q��.���SQ�Y��UА����!QH�0�WP�:�E>*�S����"g���#!�y�|�'�uu�*uA#�fF(կ�||g�ߧ��H\��ʥ~��M��3�b�*�y�.�[Y�Ң��~�
�T�8�cb�>4�:H�{i�u�_N�֙F��pq�c��Cیx�*�[P&x����A#���\��
|�P5�s@�R�#���54�I���+�픯"��� h�
i�7�s�2���!�ƌ���n�"D�L-�^^�F�N�7fʕ�E�������?K�\�8R ��P�pdG��4R8�q�V�`�Ҹ��.V�O�be��������7{�[1p�"!B�)����F�L��(.���Z�\wp���/;�>�'F&^{DT;okW,�W�2�vp�#E����׉�
��.���{�H���I[֊��B���U4
l���? XK9e�>·���PI-��M�:�Ճ2�Q8�{ ��ֳl�~�C3(������� �/��5���aw�0��J-�_��Qͬ�e�$2^�⟣�k�~Vp���awG|�k
��og#b��kBx���Vz��[��t��*�ҽ��vv��e�� ��rp���b���Ft��@%/"��e��Da5��1�XG��Wj��ޔR��͗���?'Z��?����M+ƈɃ(, �1�b"��%VXU~��yH�X��$�����4 �j9����J<R���+��Q�����x��wisп��@F@�2�y����~�r��d �Q)��A���СR['��n=��x�b�Q�`(cR-�-{7fuJ�Z�4��7��-	��ގ�(����}�����=�Q��(Ŝ?i����A0���>�������7�g2�z��v�*8�/����L���;e�=ۛ�K
�p�� �<��������8g�ˣ�T��#��;�Ba���;���l$�ی���X��S����#��Kq;�f����aA�{tb�o��yn�f76�ܐ:�o*����#릟C�*V�`��>]i��i�f���\�@yy��626¯f����ه���nqR+zHt��5�rGGkz��d�r-���M��l�/��oT�d�쇿�3�"��!c��=E4���;�t͡�,� �j{Y��o2���D�a>KzD�(թ��M4"/0:�O�_ �ɕ��P��Lu�Y+)��Y�A�C��[�`�xҨ�&}!�)�����u�}{"h����D�k'}��JO���Ca}[�����7#|g.��z���kE����.�Gᲀ^wM�}/&s�쮘��
�
�������cp��}��f(�D��~_�N5ӻ)a,}B��]�g�]iE��\^M~�xLE��h!��.��P��2��L�M#a��}�^w�Rh��*�T6 D�M���Γ%c��s}_�ƛ���$|���A���GC��l��"�d�� �;[�&1H)A��c�%ݠ/E��n�ML��v�]���ջI�^<�¹ЗK�R��u^����2D���Թ�@��٩���_�Z�3��|k�뉤B�W��W�)P:��E������/tϡ�BD72N�D�)'oOx	|�0���mO�]152J;=L���e�%��� zX��*�����0p(�?ݙ�`�7��9ߐ9W�L<���3����S�G��3�\�[�`_<ǖޯ՗���HA��U9}�"�o�D0�bG��+���y����e����	Hv P n.	s��Wނ6���J�Qu�"��v��%mkRp@��OO��1t A�Wr��+���D'P��K&����$���-�c%�ޡ��3� �����G�KqKp���m#������}$5�iL���*��L`�iқ�81��i҂l����3\���<P�i��ॎUK�Jw�[�5��ӽ6����G5&��6���^h;�X�c!��Y0O]��Z�Xl��n4�w�m��6��"�CΝ��(Wn��;���mNz��>�B�?O���\��
��ZΫS�َ�e�'��H��>�/)��d�R������R��^-���E�᫵k	��o���[k�OG������Fې�Ɯq�6ʇ�0�#�9��#��AE���=.צ�h�G���칩�������~���o����e͏%�p��R�t�V��X��5)Q��:�tYr��8,_�����Y�f��R�c	9��+�S���+���=�K�'��_���}��X/A�k���ta�HfȚ���%�-�uӃ��t�nY|�iT�ڃ���#h-@� �!��'��.
�UC�ARF{�p{�h���(�c�Cz��j ����> ��^�p��y#�~xLъ��7�a�iA��� �ȉ���2���}9~��z��O'1��G��n��k��[�t�/C{J�-�?Iu=�6I@�n�LF5��roGN��Kr�M���0��ƺ~��2��Ѥ�����@}�]�jאm�O���O�ň��D@%�\���폓j�}��q@A������� ��S��wCf6�kR?���sC@�w ����7�k�#�3P���r�r&Pkh3�a���Tl����6c3�1a��A��B2$"�p�t!�>�7�9����B\�\q���wl�!���0t�k(dԞ��>w|�{���
] �2��;e��	cJfF�}�y4��^�֦����e����^����E }��ښM��J�������Ў�2f{F���o�]ö�C;�����)/3AO��J��5"�Fw#I��d
ˡ�M5�Ě\��p���%�����{�F�L~I�'���󓟢{s��n�\5�����Vo�tU�p�<35��4���Q�������y�]�"Q�~"���l[C��S�.��S������WX� ��6B#!ۊ��i�?*������3�#����#�&�9��������`��s���*P����b�/	DqA��!�v��m�^�_�o��vd��-�O?�	�������d"=:<�#��m� �=��1nr=sU!Ћ�r3���&��M�b,��&�Ex*��P�>	��+-���զa�oF
F�8��7KH�BF����|T\⑪�6��Wf��;"�m{d�l�A�����##�$���Y���G}�@��={V�y�K�i��g�9M���}c�@578��"���T.�A��A#Zi�좞��/�H�t$h<�]}�Z"���_�C���ӶRx��$S�"t��մ2��-�`��}{fl�l�6?4�"z(���l� �Ւ{��J*��P���]�g!ƛLNc[�7'�RF~�K�);e�X�u�ۉƄ�N�et
(��j_`޳z��Z$F�L�u�3q�&�?�3�z�j�y5:УqЭ�C#�RJ����;?R��"m�~=/��AB�9I�l���ש���Tk�J�"v7(I;�uP��Q���\y_�R������'x��X�9���+�lՃq�/���R��r�~%v ��������(GLj�ERS� p;cq��|I��(6{��LA�mD*s�E~ջ:Y�@�x>>�2�X���'�Z����'��/��c�@�P��4O��9:�n�ceI�����q0� ��)M_��ڛ"48Ŧ��E�٥�˷Ft��JL�[B+2�S�U��œ2 �E��a�J�;Vb�VjݤR��X�������,̞��&f��)�q0-v�=�6OW����?Vc���oN�T�Zv'��i}8��Q�لk2}��r��W�����aѐ�,�%Z�����5䤙
x� �
�"����H�ف���>ix�h6
�NKB��WUPeq_?���6Rt6�6��m`.���"o���ĵ�
߀��	�[��5/�OP)B��j (1���=�4�%��K��\O����k}�U��6��MV���*�ŽF�����K�s��[U�[�|$P�bH�$�;m�דN0�+�s��9�ڢb�1!��җ�w�s\�資>N����
[^{��E�]�U	I�t}�\�	@B<��՘��<�jf�C��2, �u[�ˈ@�T���ْ��yE�M���ݛO�]�Iڨ6Ș(���q
��L�"�\/�?��OU��
�t3�&��K9����<Z�~X�����gR#�����QBP��{m���:C�M�����2�:I:�V�S�/y0�$�Y�5��3����1���� �b�Q�8,�0}X�|�8R\��ܵ�i+���.j�:�<��������>� <������t���;��k�C�QF��/�}�����MmA&�5&Q������\���;> ��j����W�Eչ��35z�R�Bnl�T�l|HLg�3�� ���X�sͻB�D�2��5Oi���kJ�oEO%�Q�A�W��C��L5�Ƌ� ��/���^����=���� f��Cb�|¯fb���Q��c!��^8�u�@�)W�"��Bd���m�
<��N䇗�m���'����Z��)�� �K,QP�6
�Cqg ��@5l��)_4^��^���K��u���O���>.eCt�u@�u�7f�,iۓ⒛��rd,��Ȯ��E��>���(.8b�m�g����3�� M����+��)X�Hϟ���V��[��Ӝ��[4t��Xx��`+l�'0��w�-�>�+k�_;�u��=�)6��᧢|�X��W:�3���e7׍f��boN���WFK����d�6Zm�QhH�e�B�6:\�\���="��+O|��]Kn���|�y6Ci��lM��������E�i��a;�CZ�������|��Hf�3#T���ˮ���\�ޚH%R�Ӳ��!�Pk[�Fh���	)q�1ӛ��t�;[ث���;�'����(q,wZ����ey1�m
n�`�V��5ik�4v	Q��;s�_+�f��f���ͺ��OP�b���9{1� :�W|A �3#�9��Z�.y�W.-���q�)ݘ�'���.W�0>���4�mdb_\\���ۜ�Lf����y����0[�'�Z�Zc�o����8]A��	��]����"�2�彡�����z���ē* ����:�*c�����?�KƏ���3�z�8CG6QN;�c;�<O"��,Ӯ�h"�0�&��24�+����O��/G
�>�-��[ q�� ��[w�3���t�_�c�N)��R �w�PTYA�
^׳�Z�E��@�%��:(π�}�4��5`!���3����`y�D�ҫ�����.�^"o�	bPOX����;ْl�\���о��Q�O>JՎ6��Hթ�Ȱ�p��<Pa�9����_8�vLWK��o���bv���Z���C��o�D�jlƯS�RV���V�3�f�r\	�m�ポ'�����u7
�_�X�.c�T�:�s��$�%�.�M
�%�fј�
4_/��C�����>p6E`��7��]�v�1��p�`钽�~���(FA"|)�(y��6�ɑ��.��ek��r�� �KF�!�(�
ٸ��5Aj��=��
��ӥ̶\\f1�K7�p�\v\��PC�Y�����J6�hvu������3<�m�{c8tu�'T�s�~y�۠����;.R��Z4��Q���F���GJ�t�<�˙ 7�	�,���|qX*�K�����?��Xo��g��Qxe�sUz��r�����6�L��5�E����?VC��P��sXJ�^��z_rJ�t�caI!ϴ���
����^��%���V	���0Oȥ��1��n��"����(X��Ꚛ'V��D*�*0_�e��;���1G��ʰgsg�Ǩ�T)�Xo�g��a��KMV�}�y�s^Ɛ ȠZ��x���,[������y����=
�B�ʥ��e��bk���M,�P���?T�o�00�C���μ^��F��<�����Zf+ݍcU����N�-G�Ŀ#�.z'*�L��B͔�۶���#-��M���-ߖDؙ���K���]�f�x�4��⧬��]eWFS6��T@�>F��8U^Y��%:��	��ca���̘R��gu �� ����1	�BA��7� �f�˳|�b��`ɋ�1�m�o�=��OXii�fQ&��(}�y9�_�/٣1vؗ�4�&t'=�	�PK-З��K�N����i!2�����\k���	�Es}���� �_LL�mY�bO���/��im�B�+�nAJBnVZH�%�汯�mƂ�cB��e�i�/�]���t�4Ae<�?71�)��ڙ&�vYj8���+k8�Nx�T�&<�ȄX۩����' z9�E��'GO�Isp�G�çHrŇ��<�ƗG\����ʢ�n"���XD���9|��(�5��yG��F~���kv�`׽�k�U���B�bR�W���v�u@���Y��W���֧�)?�ns��Nd9��lc�,,�d%
�J\Ȏ�.���ɮ��*c��A/��s3��O����JΫ�i6=Rt��k���г��H�W�ut�亜��g�����Tzﳑߵl���,�k� [H{\�!8ȵ��B�@��qr�8}:�Y�� 5��t�M/�M{*��xvܿͣ�{�r�v��8-�|��a�&iʰ���T�3�olH�(�RFH4(��J��NQ� ���ʖTT��:l��~G�c~��o`l~WXa��������@���*v���m:��Y�<��h��B�g�K5	�26P�T��cS� ���4���I�.�gҾ���]t�L�8n�n �ue\�	*�*"g�u$�����I�f��PF�eH�|bx�{�/DM��.�:JQ�`���̅��/�0���
s��i���%U���T��$�u�֕o6��R,�t|���]��e$Z��im]8_m|�G�D��C!7S�HF'D3h{�ԛ�j^.᜺K��㛥�/)��:\�N���)�3�V:XNe $�.f�2{K��z&�Yh�\�;\d�I�� �7��5k�^G�	~�r_�g*w�AYè]a�%�(k��(>�a<�x�E����>�a���_�����M�U�Ҵ�33�;O�x6��0q	��j��$B���q�R����V��I2"�G��?K5>�!"��z'5�i������sT
#�EnL��ܚ��D����P�&��r@��sY�"]Q!��E6��w&�0_n�l�7H/h�!L�>�$�G ��]ǫ\��x�T�����NV�O��~Sc��@��龭1쏢����9�u��]������C�ls��)�������2]�s��1-� �k�����dZ;|���������4�� BlDH]��[���`A�>��11��k��`��>��d�q�qH�5�%r���o���.�{���B��Iwˊ>�ej�w�`�L-#��M��ެ�3�K9��h|K���NY$�w�'X�	�x��q<����׍�e'��~���)+�rP��\Bn�jS{^ B����_H�'"��q��XK����4�F+��mm��q������@��ج�;��������+l��6�U�`�Ԗd�naT
C"Q�$0�����4�i��ݧ� ��h�r���E3�+��Ef�5��咝0bx�}�7�Dp�����f��JͿd5�H1i(
GqI�.��
�#���Z�[��˕!4���E����S^�|p�5D��W$|1��0k�1�?;�f��C
"+$�󥋇x��{5� CL�ep�B����C��-�r�I�E��7��Œ��,xW�F�S�N���3w��oMp�8��o�:��
��,5�~Zy�C��vS��-��@�LGA����:zj`Y��!4ӝl��%�ݗ�a�DMD��G�q�����i�Q�h�n�Yů�|L�×� �*���)[�B3Y��%Vʙ]N_��!O���$���������P=7��(���z�}�r�>B��XF,�����{����}��q�1^Wr�)?�K����e�&�n�t��E|�^�^�f�3�w$�ۼqhߙ"A�� y1m�~#��x�����j���aV����8�aqv�g����(ɩ@���iӆ����܌x��Nt�O!��E�t��R�^�ʷ���1�=3aA���}���Q>'A�ߡR��m|�hD�o�D����Tf��Xs/�VZ�K��`�*fkh �6z���k���b������D�G�M��%mH� �O $*�d�Z4�v����b�m]�\��Z��6�{@+�Mq8����'8n9D��W�HƠ�����ӛ��|��P	M��P�D��rF��W��h��.��V؝ ����d./��`�s�ܰ޶�[����XVB�C�����!0� �R�����捬�����K��eƩ˽\4��`<��{'��xH�yA�(C��8���`����3�=�:ef�U��H�s[���� y�㌆Ƿ�F���=/(fֲ�Iu�T9�y�8��g+'������e�� �[�@L8��Y�P~zo�I��{������ �'��A�^��~6!���%pƝ�{k��W*��7r?��:�~�.��W��*�JCUB��;k�X�J@�D�"0"�k�R����.�ʊ->u��$%#�����씚���x3	8�u��	����N��
Tߦ*�:<�����!�k��P��Z�t#��{�@V���4Uz!I�?9���f���2�յV�\�Ϥ�r*�xV#ln2���\�'^����6v�	�&-v},d�1d�k�Sꄅ���0���.+�m-���� �]r{ �5eL+����Ş#)���};���F���C�x�GV
�[��S�m�M�HQI�\��OJ��pA���${\� �$ ;@�q��jS���t^L
��EE<%��S����_��H��QX�ψ~����3���TOz�@����̶:��`�h����f� G�\�ș�� '�28����Ʊo��Mv��bl���K5D��  �(�cA��M�Y��1���@CˠR����a�`��Z��YE7��c&,k̾���t��~TKI�d(��0��-�;Fgp��b�_�T)�>��m�?*7|Z�m��d���[U�1,D4Frg�ug�6�Ҫ������Y����\��s8�f�k�:/A2�.W���I�J�>t���,M��T���.���D�#�#{�~ᳯ�_��ײR���ݜ\�q~T�ۄ���D��2,���Չ���HJ��}����� L�%����m��`��߰�z�Ë%5���\�rE[��a(����	��p\֍m�W�ʐ3�G��J"��}��yʚ�M�O)j�Q9�����s2�x�M|��1�j�N;{����[P��z����'�7������	��`D�m���n�ĳ���th��J3���$��G>�����/K�4��DB��]�3��Z�����ey�������>�|o���mZ&
x�K�
Ȳ�P-XfU�kmqw�[��*cx�ٳʗ���P��"vCu���O�6(ֹ�~�bS�&��.My����Bf<&>D��������A���Xh���� �;/B�\�y�\�CQحMDD&1� �=Вܢ���_��	��f_"-d��^���%l`�)���ؐa/��q��߲�tb>�"#D�Az��ڸ�K>�c^ ����xJ��a�m ��s�0{��U*?��#5�4$�V6g�?�Q-�+g��x[ �HI{�<�Ϣc֯̊5s5|�<N�\�Vz���\8!JE܃�;HxS�0��ժ)����r��A�B���AsS��]�y&�L�qw�
��c<+Yd4���o����?�#�rD���r��Q�p��id�4f�=�P���C0����B^��i@�^ �@z�@��=*ڛ$�H'T��ag�=�6±>@;>��c��i�� �&n߬V�Ga�Q1v�OZŪ�Җ~�����̤L}�bt�*NV�)1kծG�;����=_��4ƕH�	ڣq;�~�E�c�(��gq�O2�����b�T�f���"z��M���\ૻ�(e��7�Gw���_Qc�V�]�zM�m �E��k21S��x(��ޞ����H�M�r�}'(S4��Nߧ�m&�0�QX����y����Z�6�^������
y�[P�A��>������QI��ٴ��4?���u���[�(3!켣.����u��������d� N��rb�#��U��^�@�e����B���m�oqROoU?�����%;��P@���X����jw��a��V�!ŖT,��B�t屁��J�{!HH������e���#���ש9isK��a��l�WPb�CsƒR����/]P��{B9� ���ym��1r��Ye��ܹ��l��~�d����)�'oaoj�"��q3FU�n��u�R����b6�y��l��8�-�&۠â�ܢK��4K"&��s@���C�_�|�o�E���ޝ���R@�kՑ�I'���;[^	�~�|G��2�UR�=h�~�;A��U�Q����~�|��R�?�Q����ό��n����ln��S8�̠)��*��7UW$�U՞�
lHd�q�`�1�,����E�Ѫs�[.s��b�����;'��z�~P=G<���+�l��K�� ��F����C��#euw�ELOM���J�[����0 ʆW�֌�.is{�_�ϡ�g%H�q~��g4�s�樭�m��F-��ޢ�v5*��䟸=N�yzId�27�J����n��ԛL��G��C^#l�8������ĩ��i�[��R"���ɶ�=3(�g'V��e6e�����9���~/�fo-ݜ�-��G�!,�d�.�2�ו	4��#�!?7�U�hO��	x�;�����;-��>0l��X�b����ۤF��>���=x_̊)	��ϸ]{�pԱJ5�"ˡ�
��w�ɫ�,��B���A�!�i�d*�8�,���9��Ƈ�ֽ=r�g��M��A�4)d��s{<f»^�aJ*�p�1���)B�נϪH��z�g��?0�[|i`;�|�#����MY ?��W��ˤW�����6t�I`�V��S^�$��0��(;�.�nï9�G�~�Ao��JH"�wJi,�s�A��]�P8?��FR~�-4�Q/
kV�,[�%�d�Pm�i=� !S���4��35�:�E<X�����AI�54�������XT	��`;F=yM����f�O��[c�A`���1��0u��&Ad�L����F����<��n��%bO��O���aM�}�Đ�� ��e��P 90�N�*]:��o�I�8Ƽ���n������>*Olӈ�x9�w7jm��=�+N(�n�"~D�\^���=M��`����q�H�V�d80b��O^C�Δi�g��n��'R+Q�ps4.��7�`�$�7	�Ü^���-@��T��y_D1����O�1a�����=�����Y�"ȅt�bR��iSX�m0�� Z2� 5�/�Up>�շ��,i!�8 �F�G���`���V�g~,k�)�h 2�{������EP�${���m��<�rK��XQ�@�{3W#�d��o�U���ʭ�w�+����{��մL�]J̥;9��+O9�{is��W�o?��_�a�?���4Ln^r��d�r ��	�,&4�'�X�)z��X<�QxwiV0��B��3lq,�w`��M����|�zO�2ک�1w�ը�&b�������vܩ UMmk<֩�|�Ӆ*��_wm�>������^��̣��O�����4U���ɞU���C����q%���K�a>s}֌n�,�@y�ۨ��^5�Wl��+΀����Ou)�E�5�&��VV�{�?��7���[!貙�$���9�bh��b`��8H%�B�7c|����X�����=�I�O|�� T��W�8����J|xf�x����E��G����C��zQ(�{�H�!O8�>�1J�Z�ou5��w��c,�����y�\k�ݬ���b1�`�Ippo��Ǽ�-45�����ݒO��>�q/�����k+�X$��ב�r��7����my�����y>jt���a�d	����GΨ��ޕ;���v^Od ��J�O��'�گ}�\��t��ͯ����=@����el�qJ�X��2L �2�tY�6��y{�A�P:	acib# �fܔ-�dw@s�D���#	���O|prC+.�E��D]�
*R�����[�V�a�:�_�W���h��V�G���k��u:Y}vih`��W��m����c�v"�o2!j�e�sh�!�����0t�>�NԌr���<<��; ¶�i��ǌ�6���-�����.�α��.����u�C��4�p�s�d君���|G�m���QRt�����w;���c�]wAO׷���TFכS��uA��U�{��ό��1��0�-�����������)�a6*�~��#�:,�h�����u���	>�H�H�&��~ ��Ev$,5T9#/�^��<E�EW�;3ɕ"��p@�D�L�_���$�\��b$w��3�k�N� xیp����J׷��}�:+�}�������74��H;�5���)�Ea�a�ʭ-�I�*1V#���H3�����85�6í��Q���:Q@���DP��ԡ5_�{�	�(Zဥ�y�9��x��(��o�7��x�9��ͻojιU\�6��˯�*����k~�g-a������`��s�+g����u���F��A5�b�S����F���UA]�:�ձ|4�R|ն	K=S�4=_���Z@��C����5XC�`*�K$Bd��1�P
c/Z"\��#�N��mK&[�!�����ݺk&�%ĉ�9�홮yiF��k�x��3��oy���.��P��TA�}�(�4���2,V�68$�F�K���$�X���=(lw��<e$r-˂���J���a�S%BfQ)C�!5����_�5�V�2k��ז�l2�Q��檙	�/~g
��ogѺ(��f50�i�dNÔ��\�,��n'�FN�Hǐ}BZvp �r��k&�q��/;^��Ϫ�3���k�Z��%z��Ǚ.5��Q	Yϒ�*xK�TO=�lpB�CY6㞊�sd�H� I��c�m��'`r=VSv��F���)��w�wY�i�����1Ø��էD@r��H�E6�d�����a�x�,������y�*󦦼�ټ���$��wڷ���S��&u�������Lq�|e�ٍ�q���~|��i��Tq*��
����^����@m���2G����-�SRN	�@.��;`�M(-ފ�	۔�y��T���_"��|߰�*P��{_�t���ǚLp<AN�I e;�].ftŮ� ����6���a��:���6��H�G��Kl��K>V�ӪWF��cQq}�����lQT����̊�v*��C�u�J�0�+Nlz�Niμ��gx
���dȓ��x�ޞjez�UM"�+i���vI%9r��JPl6�(�3��TB.�1���Mj��S���HR*� ;E�?_}Y3mR� �xQh�c��T�M�\�눌��'�W,Y%T���ZW[�Qa)�O�]︧H���C�>�R7�S�pz1x�4�Q���?{]��7m@����,S,�W��(�u��ލw5Bb�wK��<�ⰎcKQJ����O��=��z��1�WX�5!t��*�[0�hC�uE�I=n@���$�VF~�H�V�z[�B�w��>ӧW�Ld��j� H�G����D&�r&�0��9��5	���(ihy��QxI�vB�fI�%`z�7���$_�IM��?h<��n��DD����ġ�49%�=�ݙh��h�7^����q����	p3�@�3/�l9�gŲ����ef����k�f��mq{jB9�W�^������c$6P�{@FفJѹ�y�f��4���2��3t�����pA��?�� l+��3�={�o>2O��'Vw͔�A����/,��{��쑯��In�7��yc�	��o�t�pڼ�jN�_�c�P�^�[q��ַ�I1|k��H~���*
Ǐ���k�����e^ڠ�N�Rud��V�Q|Q���c���m��RfC�Q�L&�8���a�:�P)	�8�ٮp*{hhN)���
іy�fi
�VP'���OY_��{g��/  ���Ķ�|$KF�}B��B:h0�����<���9���4&TM�[DKV��U̓)���T��L�x	����za�OV�n.�Ơ�10�J���Yj9��d���y=��3̥D�kaߵ� jt�4C���
Ñ��'mӨ��_A�s�o����Ƙ�OD��A��&K�����hM/�jO���y��*9�٤��n�Շ��H��K�3�	J�މ��d:8��<�g+��^���8��u���SF�@�B&�O9352�|�s��s�on�z*WQb�B�fĽ��7�wd��>��YΒf�8������O�+&�ո�8!�M��Q8����^A��F�\ih˂.`�����D��� ���	?�^zOqT<uo�/�W���S� (�����H����M��}S�X}[�*#�7Vg�1d�߹���[��.|�՘t�4}�)�[��{ج�?���x�����zf	��X�#���>�o~��nUgh�u�ཙG��p�p���U��_hJb�!���WҵCF�N��}�|!��oԚ�Z��'][=D����a�'�Rb,���^4�2G:֣�{K�X>	s̴4��LG��fxwgq��;��W�o�d�Puh����3����A��vb���'��q��E撨)f����Ҡ�[}j�K����<Nű�1���o٧�к�m�0�E�'pol�z�7��n�?���IKP ���$�Oo�,h���zh$F@��n�bEZDg0�����Yޱ٬=I��]a# 8c�F�=��˖�r$�7ٹ��� ���x\/���yq���D>!S��lcY�-�ד�i��#5��v��@���^O@��0�.�A5����#� �Oj%7���L�B+D2_37�� ����_�(��xoyL�t���{<כ�?W�o��*�����/�6a�nAU��An�/�#�������^�8H��('O�W�/�  6�v�fZe{A�W�� I{�:�d1yq�Kp�E�'�7�oF8���M���ח◺c��Cya��[HrP�ڥ[��
�����k�[�^�&�@�B��ț��gP6�ȍXܚI���]h6|�W���Վ�fϰ��G{x1���jeJ�F���]u�!��Us��;�A{w��~(�&�r����}}�~޷� �R����Mxt>�P�lI��ә��NG��(�OAƧ7��:�z`�1�;�/�4��������=)��T��-��G���K"W#���:j���?w�ˮ�"52�r����C���ԯ��)��87Ԟ)s�&,��$,H%H�j�Z�E𭚃��􂠰
8YWb�eb�P�#�qV|�E1� ��\G��؀��ϥ^ci#��"vG����2 �2����Ex�#�$Y����M��
)���X��s�r�,^��bp���o\��O>� &��c�*˔I���[����A��t�� D����-�TA�Y���J�Ь�Y�K�������m��̯(Ё��a�u����(����@]ϯ�����W<���sB���Q<�7B�u�n��<{΋i�Kۡ���<���"�s�i>5)2Q�]>�Ҥ���~M�	� gK8�X\~&j�_�v�w >Xɾ�v�ơ��?��N�-nԏ/*+�'f�S�uk|�u[4�ƻ�߃��ۿ	#/��m�T�f�����,Ɠ*�A�(?��l�@�����L��E�Ix�A[4���Α9|�w���: �'�ۣ�T͕�K��{՞j�Jp��e)�&�ǡ+,��d4���pj�x�ѵ���-�0�΀!Qd��Zg;�g�+$��>^�J�#�-�&`?�J�s�P5��ᦐE3�����u[����5����]��K*�C�t�V>z�7N� �M�1��6#��V���G�dF\{FUtw��2'�m�;���`b������s3����7��GPk8Y�ƯUNL�=u�ݻF�cf��x�Rf�R�5�S���J��� ڒ"ŤA��Z�@�+5ч�"����v*EB_�P�π%��~�s݂"ݖ���� ��� {����ٮI�gŢ��v�������'�4x�ÓA��w�Ajn���fG��2
�7B�d�*P?&�5!,&�S�X1��)3��5k���4����tM��:j��X���}���_��c�<u-��ˡ?��n�?��1ʐ��\g�y�d�V��?뾠�1S�|�~��b@��f��ڹ7�P��'�@��/m���7?Fۘ)n!�. �@��9-u~��X��9X�N�Cr�e4��m`i��ˣ�0mT�[O�g��'E���ť`a �"�����"h(���䍸**l�ؙ����� �^�l�nÏ�N�SR�N33lH�pf��9dPTFZ����׉�i'��$H9�v�U(�U�I�b/%���D<�9�TKݵy9&]���y�W�v;.��y�E:'��?R���r@Db9;��j� َ�k( i5�	f;p^y9��縬{<�]�EF�<�p���"�P^���jd^X�g�kV�AޞW��L��=#ʵ��O�5�\�ҟ�W�}��Im,����]9g����$6J�&.p~��G;��$�9ܮk��(���?� 3DPo�6�5�t�L�3,j�y�RVJ�y�p��!�Gh�L�8�!�˛���'s��.�w�`.�L����z��^BuF-�63��W�ۅ"z�alH6<m�pL:	�ޜ�l���>�d�ы镀t*7��6�:�'y?Ѽ�[���o!u�6���g!>����(�s͝E��d�K��+������m�e�>��pN�pd%GPcː��N��*�?Ϋf���H}CLB����_�z���֛f�Pu���q�{�?�[C.�Y\1�j�B�)����҉ �m�r!Uv�\�(�Q��b4��^0�.��ĕMNrY6|��VW��؜��`��,Ec��S��==#�1_�۸��F�+��%���|c�r��B/ʀ�����9\�Z���9%]Y�u�"�U����Z̤�
�bcD߆"I�����a�t�I��4�%�:]�p
��D�j-;^!P��n]��~���F�o�3�k��N����I;ʢ��w;7T��C�/%^�6d�73���HQ������B��Yd�F�"��k��`*�<߼�Y�\k��T�^ ^
��N6> #ͺ����vs&Ѹ$
��[;u��o�ƫ��j���.�#މ��sOJ�1�!4G��R�Ght-��.Fڳ}����'��4o�/7Րo��U�����y��������qm��P��[���������*()�\� �����a�����w���	�gI��/e��T4�w����Y5����zKgȖ0R�O�,��{ۢ���k:B����,+���V!O�)��	��紿��3b�P��m:Ӽ:�ӳU	-�~�׊�����V���2�6t��r��ku�"Aqu��F� u޷��J��#/uH��� |魛1�x��_�U�7�aL�uymr�%���!O�ߌ�܁��z���,��|���;C�l�7����}����1+յm}��d32)��"O���0S�}���]��;��?R���v�͛��Tg6e$˦���+g� �$e���[U�t�{���=��7Qp���5ګ!�f,��'�"�=�ه�Xv1h��
N'���C��45�l���o#o�2Ę��,�IT�Ud��#�<m��c�)�l!����/��q�>�\�*���<]ی�_�W�9B^=*�H��6�W	�3�����S����6��b��+:m��V�����K��������?c�$�ֶdނ�@;�K5�b%���
ȵ�>�MR+m-j��B%��;k/�@14K!4x�y
P�_^Fʠk)ǣ̏ϓO�ζ�7�%��>��g�*(fc�$[@��ۄ>�8:@�צ*5{ d��f}��Vp�Bx��(�b�8��р�e���fg#&~,��vl�w43*��V�����؛kNv��3��*AUJ|�9�c�Y���,�&n
8���`�3&�s%X��"�WK�a-��`#�eiS�親`�(h��t�7$|��c_
�q���b��_��t!3�?��	�3[Þ\dl��4Np��ؾ�Zc�a7�\_Vl;�i���~ʏg��\� V��)b2�B��Hn�]�(t��&~F����T�HN	��bs
�����*Q�k�xN�׶������^a#R:`5��^����B��)!i��&�H�-�Kw�w�Y����ٹ��Bܵ����>8�hr��].���B
�dr�2��N�R'-j�V��?��U�3*u3�9'�c�*�A�E��^n��"��;Vs8��~:&+A���p�G
_7%@ ��ZvA�T��ڱ��"�Uj�?m!p��f�vN)�rMz*��!��XY�4��i��1� �ٚ��l����k	u;��J;�<�髻SR�.ˮ+4���a�Z�a[�	�-u����{����&����4��ˏ�+�R�d��Ƨ���bL�^
�b �h(��._4���Jݔ#@Oܩ���A��weF:��5�ɰ2{lX�i�m��T����7�<������
x�� �S�3��g˄*��]����{�/QE���ȷti��X�,�CH�~�.�_�h�8�i.u&b'4r����wt�<2N3�$�KK��'XEk
�h�oEX����n7܄����F%~Q��UE]%�H�S���/�F��"y�֪ �����]I�Ȅ8W�ӰK���d�"�/эA�U�o����p���ˆZ|&��rRJ�K���(~��j>��4��Y8�(.XQ��\���M��Xx��{YS)>n#jOWIN9���jmY�.b��Cʰ�_�A�'�E��<T/�|��q��ǀwgt�����H�_�8޷Z'�LX�n���r��U��寖X����fm���&�y�*�if�!n�c���t_��Gj�=0�q��,ܢ)A��+�߳	N/��B�QG����O�d� 5�e n�A75ʗ"c��,� ��0��{�~�L,ƓxR�ݥV�CC��:z�B����k���UZ:�8^@�
�$P����⥶��G��u��FE�	p*,l�+"���5����t���7�Xv�?��xk{�c��_��e7��>�S �u!
tMpHv��RӅ���(k��662��7�F��^����_a>`���uR�8���4<�;4��~��uB���EJ���/g�R��T�� F��v��;��%' .u�X7��=���P��k�
�ʭdJ�(��	�4<�>�@�Bn�:���G,����	q6�)��Y%�XPD�����C���웝~�W�����^��*P�g���6*��:�W2s>�d�k���)�Wp�;��!�.�|f$A����W��Up��qa��~+�|'8�Wa��טA@�1��Ĥp�8/c�ۘ���2�+��kВ�q��=�)�yc�U.ju�z#A��_2q�y�|�T�x����<°�#r����
,�IC��iF��[v68b�R���|�,;��)�;Q��G�r~�I��g��������G3�U|<��D��g~���[��x�H�zx�0�Ԭ���0�ﶢ���0X�uZW]�c'+Ik�G�]�V>l������~���I�7��j��_��W�xX�����W����J�Z�Tx���4B�5kp����Ȣ܌�rp������k��&�]��z��D����}Zbѵ]�U���"m_�N�s0�g����"Վ���ET�� ;α����������z2W�v접���H���:Fa��j"����C���h�ӃLZ��	w�`��m�p:)����dHN����!vi+�� �]ۋ۝�L�����Nm�T�U�ī\� ��ja������7sQ5���a`O��]�@~J����O��M#L���s1.���TQA^�;�ٮ"|��Z�E����� u}�&2�!��A ���r�� {=����Ȑ�ݘJ��WqQz�2�|�&�7޸v5��u�Z���?i�ŊjfS^�Ƿ��y��l������&7Y�j��ǒB,H��6 �x�ʵ�Y�):f�/:�GlL�}�m�D�ji��a4=�5F���}k����c~|Zm�Kn�H���c��$o�4A�S��Ժ�����?��h�s d�hjh����^:(y�p8� ��f����� ٬���}WKx�[4�%K��x��Laj,Q��λ�14ﺲ$��*��I�
{�{<B�u]�"�l�$�4*ђX昍d�ç��J���I]p�TA��zBZ��m�x(	u����l�پ��c�1w��|��� ��	���z�!�$���s;W�(��\������w�:bmU����ǀ<�k�w�g  .��A�~~�F�p�`�C�mC�ꖱ��r}���8i؞��<�����	o�� l���9�.�������T@CY�k�eBYl�!���:u���ʔ���	,�T���ϵH[���kZ>˛87�6�h��V�rM�@ٶ��C�ʯ�ð��7���y��&�s(iK�R�$Q��Vی>-��n���2�z��h�������m1ꀃj�=t�N.�M|K� �q�X%�	�����$�?b�ƭ_�m��V��_����p�O���h�dEP����0beL�X�ۤU�σZ�p�V�\����L5�h�X-�]��w�iK�� ]�$�ܱ��ᦅ��W��XN�uS�,&=��ڏ5����^�-��hչ�!![�
�)�E\���눆�ʍ9}���kf��PM@=�mp��cHR�Q���g�����jx�&4��s�W��p�H�'����� <V%��}9��M�̷�/�����I�q����V�A	���#��e���5`�JJ���S�>bS����֕�-��-��6.W��O0�B��R���E�V�&NfS�Α��Px��Jp'�ʽ�Jj�x5,�epP��R�ױߏ���sak����X!ק�\3y.nj��ըx�/��n^v��W��Ϣcǉށ��I�Y����Xs��d=?���'�����&]�	;?�m�7W��D���G�$��R��!p�����Rj�U��:bO���l���^��	��mq�o�Lxzoqˊ�� �%���F���|
����R��c�MYT��1�ڡ�E���'H��M�c f�ۧ�O��H�wg�!r!�,��U�@7__�U�B\�HE���Z�:{�>�3a:�³��,$�6�g��{��	�F�C,g@��D�IPث���8��wF_?���: %n?YtU7��P~K!�����s�H�v�Q�.����k
��&z?e6���?~�~�-$IyD9�U�kO�+��zg��.���*�Ǎv�mV����aD��u�����qTT�e*Ĉʡ�u5X�RF"tv�If��i��֥-b�.��FP�+Qu�m��m�i��j�����.R�{�n��\����d]�L��>��7C�H�q������_yY,�ʺ�n�-A�r;bs�%ĝli'�-8�y��˗Ua����b\CgpȂ�~5k���-�e���O5���ҥ|�e����s4l�CB,Cm(���U%K�̴���R���z<������聝u��ԡe�?Mw�6��:���p�J��!���SO�m��nX&3ʣ�3
2�U����0�3�$�@��!;O�AnWK�����w�D6^���������F�4�)I9�S��K5��5ѧ��	1d�����x��swo�_;0�V�-��>׊��Ki�q��8
;7��hQ�_F�N{�P��p�TYX�C�v�Tp%���������� �Usq���~�:u�­1rw��*�S!�-$f�8�N��X�1h:�.���	m�����=�^ns�g���=���3���r�W�gj�`�9v'�~|d�<���g|l������-�b�!BM�T���$�zm�p�J�L2�iR�v�߫d
����ØTxy�;��$��[��>֒9�M�?z�����/ڿ;�TK�ؤ�����7�A�Y��u�Lir��k����Ϲ���X���U-^t���O#�&50;Tg��%�sXmu��l��"1��7�T$��e���.��E��+��=�C�b��3�G�5\3y�{j� �X�o$��$� �GV��$IUݜQI��3b�0Y��6���M��EA~�^3&)�z|؀�Ye,}iC~9�BBȎ���-��Z��6S�:Լ��̌�'H��8��|2n�}`�B�gJGBR��\��	u9�~9��w��L��"k�K�&� [4*Lmc���R3ढ़���_�M�_~"g!�Tl��pن�x�hi�7��ǼX�,���B13����^S�9��]71�,
і��ɑi$��C�ʡ�7�Vy�!���~W��_�ў#H==����`�JA!C�'�Ώ��>-�(Ұ���%n)�@�ؓ��m��P�G�쨁�o�ht����}��ag���h;tX�A*�ʑ����)'ϓ19�3~NE��@~_�'�8q�O��_�k0�8���������Q^4T����%�qF�mÀ�R�=��3��q��E��q�>��c�-��j;!Bhp�-jM,��Ӎ\bF͍em3d�G�+�l`��sɱP �Ǌ`�	�ԁ3P�7*a�v�J��}%��gH� ��ns�+����/��#�t�2>D�DZQ�mB)�v�3�իG�'o��di!_� B���Ѓ�OG)ԏ����<��`L"�����4K]�� ��
^��p���54�K@�&g�Җ��V��0��R��H���x˂�ϥ\^�*I5Lrt$1ϼ �H��J.�A��ű���Y�`����<�g�x�i���2P9@�#>�\/�'0�qF�Nm��~�� JĂ��M��p#q
��_�t�����u��8>��$�[_��:X�b�#�"��8��T�lQr�b�P?��1
���8���]r:Z��x���*�R��GW��I��a�;&"l��!��������JN�v�ٰ����#I�f����f�#r6�ϵ��F�	��8��6xLL�a��%]��kC�o.�5V�#�W)j���f���]ƐTS���p�$md@O�\�>pF0Ron�9�WGw\N墙��Q�ҡ��X����M`l"�*;��'�h�@��p���콄$���W��u/ (1]qi�����'�/@%bj8	}~e�!� 
�ш?]�RH�iAY�؉������;���%`�"�^!�k���[C�y�\ݺ���]8�M�������M�j��-���q���2��#��ݘ(��V&�^��TU������>@௲=��  e�0Qu�׊cMI&z��� �=	>�q�;�ҭ�C�#tM���t�m��õ��>����l����?1J��ׁ#�v�(^���.Cq�!��6�!?���9�K�l����	��E6�+�J����e%�1H�y�S~h��T�;6&�������_j5@��Sc/k��iY��<Beѷ�����qE�OYiM�,�L��B�<wd���3c���5�%X�:�YW���q��}PB�<h�A�$5y�L���c��%���Eĩ������D�[�?���6Er��B�R f��Ŀ�"��V����oB�i'���jg��\Ml�%ڜ#��r�V:�E��9~��;*\���L���S���w*�ɐ�@]%hWU�Ą�R�t��8 Х���*_��9%���`य़��bXwe0�hN�T_�rЉ���tM.�������S�ӊ���������j!�
�n�Oc�GǑ��#�0��hBaݤ��b��Uh�B=����E��g��������HEC���_���e�`�<fӁ��ȑ��&�_�UM�7�E��,s�bi"Q}����Y"������ZL'<ܪ�R�>aR�ӻ����nU�;�-^�q�x���:dv�Y�%Mh��@�J��EF��e!g�*W2��6����7�pBv�,u-B�IE��7f�o	�)-��b�tFT`8.e7Wo��C�"s����9�w��{M��㱕T�����8]=v&�4�Ы��\�}�ָ�H�(��J�ֳS�B���&����q��Wk�(Vw	_�o��zP����u7� ��Օhl�>� ��	�⠍kQ[�x����M6V
]�m����"��D�L×f�@i��%w�zB���Dx��Hw��IIIŽ��<ݡ2����b�p�b/����$S\jd�C�e�Ŷ���ц��e1����fō��K@��97����<���D���vVg(�m�w���|�C����H�<���{sƽ�ӣ��fK�,毝i���0����Y��<�:� �VϓH�2�ҹ�Ȕ�izh���^K�����?+hl���&��UYg?�J�'��{PCÀ�7���y9�n~6�KZ
V]��,�O�s��-O��k_�br_�E��4�<����bm!ҙ�E�ɬ���gW5�f_��?�lʭ&�4���(;[��q����Tx�ȫ�'��^��5ӂU�����փ��'<�엦L�Fa���,߼�"��Ez����&�6�����N"�������1��`�q��a�a�'(s�q�܏���<l�aA%*�o\��f�M�7$�~���;�z�R]r[��U@��:4SG�����9�����'�j��1�p��pw8���sT������ujѽ�`�a	��O<�d�����_���z�d�� u���6_�6��c~��IV��^'m���ԡ�D���=��ewKy|s����N��J� �nĔ��Q��;m���`�}8���6\S��CRD]�ڮ4X���P\O��VX]� �\�q�*@.62��*�K$}�;��p�j�q(��]yɿ�2�^��/+�T�)k����zd��0��ڀF��Qk�~���|�6Ɖ �2�	Dqx;�
'B�$�.��J�nC���	`��]׉ԯx�K�A�R9O�;�?A�������&2���4�O�&��bC�M��Һ���آ�'���4��O�*,4���8ɞO��k/��⭁J,^A��[�
&uB��u�o�K��m��� 5��<2�\�=��/	�ףz�]'�cғ_�u���NL/�{o��LFs�	I�rִ���w���b�b�����ӑ���xʓ�k�QI�d�S����ɂp�@�I���Z�� iA�ݕrz�o��K�+l�G"��=j>���%K�.(�0�ǭ
��?����u��Z�"K����8�-/���'L
��Iwz�c�������'�˙�PS|E�ۓ-)<} ����rXYm!�=��i)��Ta�t{��|:���O��o�	�Y3��|��sd����|�>��F��p>���+q���w}:�P	��wA���$&q� �����M�I3�3͌�����7�jռ�:�O�bc���q��I�4a\�L9�=�G@�G��<�����sⰴ^����]CSpM����0�m|����a�`�-)(7h� ���_ �Uߖ�9����m%�Nzi0��>��3͏�7����D��\!�P����;����rf�Q�^)R������[��鐢-*=�5]Mq	�7�#�>:���eo�C#o,�:�D�p:��#_4��Nrӳa�+n���O��Ļu�j�̚����C~7�t�U����
���Ѿb�=�����6�	�h�����Z�^i�_Q0n8!��z6����}����@Һڊ�k&D���<��lj8H��v�E
���F�yN���{r��S�sX!�(a���N�3�⥞�X��d�hCH�x�̼ɂV���I��c�GJ��H�mU�����׆�C6�g͎	,���qA���$ǝzw�ft\܌`�QG��f~`5)�~�~�Ql�,����By�/�*���&�#�G#���i^nx>�[��\�'A�2�l���,��n������(X�!L����&~Ew�4�m�C��;�(Q�Þ���.���Q6�9���õ����#<��5C;�L�$ @�IS�C"�Լ�3�/'2�L��ں���a�#(yoyy��5NInx�&&�m��wf��T�n�&4��g�Be4wl���;�c�h=��ȖW�͚�x(���Ƴhա@	�nԏeO���0{�j�e�v� ��	�M[�$����?��W"��M�le�������9�av���S���|R�L�ƫ4�C���*['|言��Ȗ��ꚥ��m2�6�R�-\
 �h��4��� ����A���I�J��Ё���o��jC�f ����PZ�X��
���ߒM֫^Qv��)�M�A�)W��K�_���JX����(q�W#�����%��M@�:��t��	N�Ei!I55�_�$�J�
�A3Sk�[�4.���Z�CP�֪=����$᥻��N; ��꿱%�Dǁ�&�����H��;�J'�f�8�۱�L����C�vd!J��!�+Rj�jN�W��� ��3��|�*�<�@j��6�j����FR�E�LP	�/���{�Ċ�e1S�៧~�� "1�e�
��Y�6�Z'�7:tfv?�>bl�WwTi�=H�~��dN�L��&mU����am���q�|�Z�0�|p��,�t{�������v�4E�	�H���D���]{�#!��Q6���i��`��:�d�E/�� � s3&�� Ӡ�#���}�Y�Q�[�TV|ǚ(���Wșj����%P�^ UD:��Ӯq2f,���l�SE���\K���A��9��0��c\( .�	�����`p
����Ջ�$�@E�2.\U;3Y��^<t�6j��hsl��zvh���3�r�!��.��E��ih^�Z 0{�o�>���t��'�vr��<��I����5dk�ف�I�)��9�(���]�8�(��Qގ^Y-�pp
Ҵíd1A
���B_ԏ�G
�����g���X�D���Ylܓ�#V�>���{�S|���@��͡�J����h�>���[?$~�0��C���l�^Li~=3|��C^��?�����ź�u��ә]�_KY�\�# {�t=HPT믲��" 2
-%0�	K�����V����zO)��Ӵ��X	^[�#��By�6�H�}?t�����k?�{P��~����I����:DAwC�o 5^\8]��ךA��M�]�)�s�i�;3�	��	W�+�s�9���-JA���5#1��I�췾w�y߿��V�D�������`
�L��=s�6��ew&�Pto�<Ȃ@����Ő�^s2���1K��t��8w��o�@,�h:�y_B �|ۙ�1d<:��ؽ~BNaYN�k<x�ޅX#@(����n`t��ۺ/���zH��dr��q�4+R���AV�y<pQr��c �n�O6�-�e�ӯ#�,�V)-���BoȻ��� n���e>������}Ga�b'ȰcZ�����i��#zP���^+���9�T�$�H�����[OQ݇���k�Z� �zV�o��9�����Z��%im�ʆ<m"]^��T���K��Э^Q�鹥䨇����_� ��W2�^�J4��t����_��@�)$�7��)~�`�[���M�u}�%�k����8Z//�q��.w[:�S�Q�E��cq3� /���ȟ���H*x�v��F�ЅI�>W×�d�FwW��8�a�{@���4��z��k�E#�X��������G������0o��8��A,p������ᬲ�lh��H���K�O� S>F���^��+�W�0����&�Z�ē�+-Kg�8���	����ĖR�T&�q��&��/�P�oU������1�����D�5�Y\�onW-��ІeInÃ���5�7[��?Կ־�F��z��Ӂ� h'͡��IÄV�?Ŕ�`t���=��1{Q����ő���n�'`��)m~�7cVS�6E�N������%��u�_���
���j�@���낾�-���2]`^�����&�K�:�_ �ZMg�6�~]�k?h �� ��q���i�U������p!Y�E�_�eC���u!��$�B�,�&��YfjNU��t�X�-|C2�DE۟>�f�9|��*���A����J@{FLc+�+���7k��Kr啋%�w���+�.dNjw�ϐfs�_�$��&ޛ,ـ��B���(8�d	���X��#�R���� $)�B��Ywцq�?,��Ů�-8�	��'��z�Q�!����CuQ/�^c�Z�`S;�aL�@q�>-��f����5�^9] �kt%z.�QĴ�/�� �,�}�m6�WE.�h2v��۬HQm�ջ��[���~H�	�Sι�Ih��@�a򭿺0�X��!�4��|�%�5�7�UQ��Z�,�D�\��\ԋ�?�I�(j��!�:`��8�t�!�{�Ԗ��XKH���/�6�"��c�_�τ�:��5��H� ��$��:��#$p��KU�Ѭ�6��
��%9OC,#�����4� l�(R}'�͢�"���s�����:��a�y��)*C��$m'J� �����8�(+>F�|�Ӭ���iV��-�#�~�X8��h�OY���%�b�:�4��H·1���p2M��B�Ǆ��!��
���B�,C�5���f�\pY#���������V%GWbk�~���� ��m���O7�u�Ap��B����;�T��i���̚Z�x��j�� &�`y��5�,����N��+��Ҁ۵T�f��!|,u�.W3e.G*ǅUH٣p��%R����?d��M˻"�����$Wy�W�[:;�̛��b�0�71ZJѕ��RM�G���F��L�#�q�1f	�"�e��%8���(sEXǱ3]��#p����0����w�q�,�F�b2Ξ=f�]?W�����'+���j0I�Zs��h@��h�+�$�a�����J�NΌt��#Ҍ	'�/A]�!8�M��[��3(�I���-�<���!�%�:!)[�A������v}���7���r�_�@%۱&)�߱D��YPk�2�v��b�\�&�\#�g�� ��Ff��M�%{�E��5�nNmG"��2Tdm���k�	����ޘV.]\h��Xl�󠖾TE����eGs_̟|��PȪ�w����$��_�VfY���*I��VFXv�O����� 	�A��}%:U%m�ʗf����̣���ɡ�N��T��i1���h��RDX�W��	�f'q�zx]��{*��y��fM�٥����T-��364�)�0Yӯs�Nb��ߴ$Z�{e����E J�'n���/yה�Պmqbb����6��.���Ol��㬞Î�3�1FC��,G�-�V���g�TF�ۊ#I��m6o���]Yg��1<��k��ۊS \��]\R�z��#�R��x����v#��9#�(~D�n�} �
�+Y-	3Y�y�?��(��<��TQ�W����F�OÐ�o{6�/X�0��ٌ@dN�[�n��#fL-T�����w6�|��I��|��Q�ˑASz�&�#�ʠQ����Pӟ^OPj���׺�'3�\��P\��Z`�u>�@5; ����l<������z-�N�<����2��A��j��q  7Xಁ �_��e�W?ѹ�yW�u�K����(�x��ʂ�����y#I>���@�0����b�S|�Uo�E3d��TU�~���������|'�+��7*H@�����;�{�"���&;��7gp%R��.��M:�q�Gϓ����:�O�������u��m[�O+��>ڔ���	#)�ų! �9ݴ��xe2��o;���P3>�I��.�%39][�V�
����i��ۇ�z� G�*��4q���7�8��=C�+h�s����q�hM-�������'�%�0a�4u¡qȈ��˔�j5�bn�i����~��f���N�!��y�j,P�#Y�X��-�9�C^&�����To�����V�[J��R�L��ה5G��J*C^�_���R�g,�Ri��*�H�7�v�r×��7�_s�Y"������ui5!���99�v.��&��0C��D&��%s��TᚾUe���,�J�,Z<�+$�%毁)o�������@nh�>R#���˯h�Y�w��|��l�+��я�)�� 5�JY*
�R�K܎�w����4���|�4<���|�_}Z߰�bDX�-ZB�;S乁����t����I�S&7�V�*���`�F����!�������0Kѣewg�P�`a)�����SF#��4MkY>N�s;�;t%|��D�_�e:�-�[Q�V!��3�_YB�6��Mz{��#��
|�+�m�=:4�!a���`� E�����캂�w��}��IW�qY���L��Թ;pԣ����4о�li˕��L���d�`u�r�,�g���~������T$P���Su�7�Z�t����L���LU�|w��!ݓ���Ɣ�[�x�,�G�'-�{Ū)��5}����1��d�׹�n<�^�1�m��Kw�VKOE� �vv9R~]B΋C�
�"(�.�� �6�2 �����h����h���ozNЀ�I��#|&I�i�x�m*˹���pŧO-�9���i6|CO�'�"�H�^�jO���8�:�M��0����^u=B
�� ޫH_�eSy�Qd��Y�)=
d�$����DP��0�a,�@vx[@����s���vE<����o0�-L��[E�şa�8Z������ӝ��x�R��� �gy_aY���d��\��֒�O?���.���op�X�k���ڒ�����
Q
���r��~�uDr�5Q;�l�9�E\~f�n=C2��^@?�@3�8�e����jE��I&�p�h��'3��5)���)��$&�u�T�3E��+|6&G��zu��F^x?R�P%z���]J+8�U (��(-Ӌk��w-�V'q߄�yn�j\WKx��2���^:뚼?EVj�L��h��Q�9����4uo�ޡ���R�s&Wo5�[S�
�0��p�ߌ��Ÿu���t^ͅ�`���'�SJaӔ�4�|�#�\�����:��֫�P��P��#y+��:�g�6��pl�y��$=�	I\���Bx�W]W����9B�,,C�C*�-���5�0�`��mv$*K�� Ĩ�4a�w�$�WC����1#P�[�t��C������3�ǎhƞ'6�� o��G�&�>��A�N8�z�m��H+��h�r|����kZVMJ�Q��o@��~�N��E���B%|0[�L �<u�c�I�M Ju�
�m��-]���'b��t�5iF�9	��+4I٦�Jv��x��x�ǆօ�d5�b���9&l���0�?�Q(�y��`��"mm�K��ح��U\g��и�Z+��{>�D��NiY�0+�o�;����횙�&��. S���~�$]�����=�~����]V��q�<�#�'VX�M8�Ac?����Ui���)��Zc�V���jݸ5,�X�����N�LB�X�r��<�h�$VVτ�XDi�ig���0*�:�8��&,�%���o�*�&��v�v�ܤ]�vL%u��a���E�0K�BCnT8"�`�������W?�c�q&	"Vd���R)&.b �;�m5FB���6��;�"���H�o������n/�Y�ls��#�U�p��߭��a�Kۯ���ؾ^�,f(�9�({����C*q�3찕>b{��^:r���o�Yk�g����:�n��o��]}�	(<f		�Z0q[6$�-VL8P�$cR-|��/��Rg#ߖ�P2p������h�E@A/eYP\��TL�%@S�J�(3'�c����vٷ��7�ȓS:Y
�W��v�F�~�'j�>�%sz�4��UFj7��.�#	�t���5���b�ߐ�Ǉ��`�0��`@���&��c.���WG_ϯ�������pJ8���`4��fV�	�,�T�A�_������؅r�j���',��v�AQ�����!�~�Q��V���Ū#-�A����\y8���ьY%.&ϗ��"Mb=)��7��yJ�n����@���)��=���u%�q�Ȓ��/��S�И�|Y��gqqN/���HF^v��ӣ8.w�X�a<�Q�)/i(�[���4��R��-j�c��3��յ�kk�,���+�m�^\$�<MY̹�w&"������g��/�>�y���V��f9���!gJ�iX6_[ɍ�DUJ�pC�9L��<о���!�mȯ���Fv���ALh8�C�d�8=��		� �'�`Bj�~E�K~ګ?jXIA�BU�ɜ��6���e�y��K�Q��@	T��X�a�,*�]	q�I�z��H ��Ke�����[���x���������M7�GD�:�~A��I���3��|�����ռL�Б�OLd��\��~�2�Q��
�|���*���9�d�D�?{h6�ٛ�2>��"<��L-)j3�
��<*�\��U���n��Jh}�2�vۢRr&�Ekya:r��T�82��Q�<��?�9�8�5��
稙�3��6��<Yo�����x���Z��ȶ��N��ޖ����+��7p8-��. %�RљW.I���ڱ��^����P�j�I�Anҍ���q�\�˿��%˫�v����%I�<C�����������1F�
� �Ӛ$mF��_P<� v�ֵx�U��:�x�0";�P���#w�<*ꁳ��'�<`��ˑ�����vP��,I����i���l@Óp t�/dMi�ij`�<;_5d�Q\磟ɱ��p��%��d�m�.���c-TrB<��l'�*���k(
�1�{��
������� �ʵ�%��L���N�ٮ�f�ZEUF�j�l8�|ɪ�C2o�p	��C��Q�C��Us3�5k���?kζx���R3��- ��w��l�JB>�'�i�2Ə�h�|f^<����R�>��z�D��NH��IC�q���`_o�q�º�}0v!.\��}�D9a��!�7.8���h7��Hz�n���?�w�y�W�7y�S��G��][BS�r��n1�&��`]M�q�U���L�h����Y%���(���zgm���z��ꯙ�r��lV��P]�K�hO�h�$>�<�qu�0<\�
�ݑ���+��eر��No6Ć�Z�Q^��~�8%��._C���xX�ӷ�a�x���F�!����^&�N�sO�_�"��K9���ٰo*���jq���$���i��@�2�ݬ�{��� ȥe|1ad)���9!3{1��̬��)�s�%:Ӏ����i�:lہ8 � �cg	�W)倛a�E�j�����}�������4(	E��r�A�^�Ȥ�p�?���g��mT�C�~M�v��e�Ф�h�_��v;��Y@���U9N$���!:�k��ڟs��Ұ���#��+��1�ʇ㒼��]���b�!��MI������B%KJ!O���^U[X ��4쇲!h��m�^"�#��B����ǫ�z��HGF�k:� ����c`t
GN��y��n����Oߥ�04U)�/���7��{[% csU ԍ��I�)������ط���8�5���U:�_a�9g��%�p��|܄4�i4Y_(H/&�s.I)�sK�	�����C�יD�1[��Z&p��p���;�C����_�6��i������8�~��Hq z�`¡-*#�!�Շӝ&F��� cI���M�� �W3X�wn"D9L�S!��\m�a� V���*��ݷ���Ѝ��$�SB�w��kv��E`�}r~S<c�5984�"�W+���#/oO��t)�_�������j����?��i����;f��3Jh�4��	��j"�&;$���?63ym�PN��!�$qY�-���ْ#a���� V�?��2�혯(��:����{�^��3�9�*�2.=\ߘdj.yL誹Ӆ$1�m�╗��o��P�T2rK	������]c��+&�����b
f��^6�͊El�:� �x�1>���l��룝p�t20�ъ�8�e!_܆��|��`𫛨a^m�(��þX�;}5KUK��2cu��/�'3�t~G��x�һ%qfԪZ�����0^_a�*[J���U~^&5�߇�)�����h䇦U��t2(��ԢY�2Ѱ�E��-�إ��q��MݮdK��|�;���p�ߨ���x�R����8���u+�)'�ɗ^�b��e���G�-� �x̺(@/�,��q�,3\�owR�� d* ���CY��޶�<ݩ�.yzU9@u"#Q+�v�	�A�Y�u����n?��e"���(�K�%,Mn�^HhX��j]�A�?W*�i�����[���O_�\�{��AK���A}�ʶ?����t�n��@�L�è#�������$-���GFop��vI[��ʦղ��G��`H~�Y�R����-;A�!Lΰ7�k��Kܶ��>�M�%ϟ"��R�'�I!O�q�P���Di�>��Y�K\N�k�mQ	'��l��u^u�q��f��d����>;��Nu��6�{�`a5�0�lK�[��l8N�i�1x:�>/������EG�-�&uvI�D.	�ڼ]Ҧ�=�is6�'�9g&PtM���z����C�	�_i�6�U���1��W�
i�(6���..�2bG��^MN�yP�]P�66�Q9ɩ7��w� ��Ʉ9\�C�?��b���v�/��K�.9�@en�OzS�-T,ef �Z�T�ԋ>���J��1����Mط1O��[��V�Ҿ�a��d� {,֚�$I�	0������b6;7�i
�W�C�����JR������K3�'�^�K��v���>.�/|�dș*B ��)u%����@D��g�� �a>v·�*L`�����x�-���l�t���>
w�s�i4�%�.`�ʗC�+I�?Ѳ�� G�;H�QG]����FL:����oٽF�Z!��'���ûy�J�#Z�c�����\!�Yjj�g�5IK�} v��E�����h�ؤ�mT�i
��&���mm?�2�0��`9#�(���r��ÿ��ߖ^��"]��|F�eP�ٞ��V7�㤖;�K��3�P���lW�5ta�$͵bO��9=�03%֔�c�<-Ϳ���S5�O�mT�4� �Q,"82�� W�k̕��$"� ��-5+�@i��B�q����D��n�3'e��0�,�}����z2>�]{pg��?��5��+�m~��6��(<�z�I�Z�]M��V�Y��o+�1UVD�f�ٜg��~F�V��|H��%����T�}�_�	���6�����L�'uI���� H��_�S/�Y�A�!9����#�ټ���t�6;gQՏ�ڗ{�݆�/��jPBI�-̀h��XA���/f�m[�o��'�^Thf'�ID��Ć�MQu�o��Z_=�}�w�dt���`����&r����ie���;@����V�mxn�V�3���'>�@���Wƣ�D��:_t� a����� 8���j3���5�C��m��go���]��aԇr<����rڙ葰����^⟎m9tK�Q�˒Jw��Q:|���R�p�zx�����)����<~*�K� �l�� -��%�؉�\hN}��E%�C����8����Aw�Eu�� ��HV,(bn���Xp\���f-�fi�(K㊂(X�����Յ��:A�q�vۧ)/Ӵ��X c�(�Q�h~�gm����d�FN�Z>mϢn���N_�u�E�)���Y��я�u�l�w�B�5���+rI`A诖sG��X:�\�?u�;��a�S4�c��l���}0Jl̫�V�R���UoO\8�b?�O��؏>]�^��հ<��b�üѶ�|w��`Ћ��9u�<A�8��G�̣D6�	9�ڣ���<_����)�󙃴s��N���Cs�ӿu�Qho.�&���o� L�(�h��Ja�p��تռ*�Q�E�� 5��h��2�]��H���fj�K����ƭo�1�A�u�-��x�2B�t@�I�}$MWK���:.���G�6%��*��4ǂD�0���;O��jBC�$�����A���Q��O�	?Ѫ�_M��\�a�:;'Ua�f������9��{*��Y����]õ�i�2D��gyu�Rߕi4~��l=[Q�����>�y�U���nB� E��������U)ȅ��|���5����RЊ�JU��To�:�9������|m�Sr��aH�� ���9qM�&����X�G��g4[�5
ഉ��r.op�5�B��,�9�'U���"��b��[���߻���/��f�=B�����0��
N���V~G�S���_YM�EĘ>T_f֫�-.���5М�O���&�j_�'�{l3T����ݔj`�X=*���"=��.�Cqe�/̽����{�,���f���[� �-�ޫ#�^/x�(ֶ/��M��A�X�6�(����F�ׂ�h6�Iere��l�����2�b�v���@�?�����La���t��ci,���a�P�����'�Zw��+�R� z�xD�!�շ������BE�5˘2�"�2���0��>�eK������E�oe;+v�6�)���
�}������R����'�CT���h�dN�A�
I.��{e"�q��^;?y�.��d,����c#R$�Pb/�$[��6FTA�ϒ���,��%��ƛ/�x�������R��;`7�i2�U�ҏ�~䦳����×S'0��R�	�x!�J$��W�xN���V�� �%z����-��Y�ͿU��Gal���e�Zr����n{UVz��`;�!4??0P���׹2ZI�6��-�v�U�*l`)�9�m�C�R���ZA��iF���$���	K���v�����)��